PK   *��VX�EfO  X�    cirkitFile.json��$�q&�*B	�W���/q����!@I��� ������S]-RK���e�3�{Vewe\-�>��IJ��N�/��0���������>����������ﾣx����C��o��ݏ�?��N�����������l�������Cӷ�SǢ��5���	��LS��)���ѶC�ړ=ٻ�~����$F�'s�"ؓs�"ؓs�"�Ss�"�Ss�"�S!� E��R�A�`O�����j1)B�QrC)�H, �Rn+In,����\�!��C$r�)�H,�FS�X�ͦ"��f�+@��Ï��O'W�Ua+ol�E����b��QVmS4ɏ@nt��z��0<����>��Ǉ�����2���>�܄;+y%N�N���;=��> ���r���C�X�]�"���1Db!wb��B�:��E%����jy|�$��r_⤾�A}���/�%$�%^�K�ȗ�ԗx�/�r_"�H, �6r_��D�X�}�"���1Db!�%b��B�~#�H,�+8b{
�%1Db!_�C$N葃C�An����!� �T�A�Z3 .�JҐ�1Db!�b��B������!�?C�S��1Db!�b��BK�!�C$�XZ�X vA�3�m�"���N1Db!��b��Bn;��T�m�"���N1Db!��[�:���24R0��i�>�ۡ)�2�ۅ<,��B&�Y29H6y���b�19H�ynND����I5�^�J.�����L:R��r"&)�f9��a����A��YN�䰺�����[eE\�{��q@�>�u�}�VU���{���nW��Z��>��N��PmRU�Ry�X�����:#_�`0
�$)pj�]��%$��b�Y9�e�Z��� �r?���i�
���v2�CRV��n��q����Y��}"@�*�7�Jٸ,�!�Z��:�4v������KQ��}Dd�U �V���}���O$�*W����4ׄ!����� �`pV_x���^��e���ќ�D�v]�"f�Mq�5�5@�ќ�N�����యʎ����ce籲��#,;;݆ �!deGXv����X�A���=X�X�A���=�XٕX�A����������#,;;���!deGXvyg��,?�˻�`��t���}��gX~�w��<]8�����t�[,*p���7R��;Kn~�T
s��F�&�8ǡY�eΐ��&�8G"p���G`~�� ,?p���G`~�$D~�l	��;D~��dq��&5���k�x�%pp�������Z�����������{:�Mp����:�6a��_�Z �����G`~��A���w���o^�ă���`�]�QA�N_���o�"N.O�%et �g?X~�z3$�<�q���x�kq8����ˏ��r�@��������΅`���,?��=��CW�����ُg?��`��_�s	�8���#0�ܡ,?p���G`~��(X~��ˏ��rWT��������~�`���ݰ��/w���/��,?��=t���X~�7o�+[.N�������px�ӗ N_����^5)���a�˜����zD��~8���#0�܏,?p���G`~��6X~��ˏ��rp����������`���,?��}ױ���ˏ��r�x��������^�`���,?��]����/X~�� ���`��_>,?totsp���G�X~�O� ��`��_>G,?p���G`~���������K��+������SW���5�>�M(;p.�|ֹ��acW�'�8 R�2ǀ�:������`Q�Zy�ok(cƛܳ����8�Ό��!�(��$��e6{0fR��^��mr����g���q8��.B�C�ʎ�w�{vVv����'��˰��B�ܥ��p�C��vr�x�ʎ�j�=?+;(;~���p�A��vr���ʎ�Zu��_���\B����8B�3vѯ~z�$�fhZ��y��,�-Co�����@�P�Q�`���#,�-Co8�"�Y
r���r?�}�mC��/��α����d��8S��;о���7�ӵ�.[��-v��� ��[���L���\��f�}�t ⇦�����t�/8���;���}+xa�<a����>�,?p��w��'��[���;K�%p���yD~����@��� �g?X~��xڰ�D�(Lޱ�w�y(�,dd��dkz�r	��',��Go�h���\q�s/v�R����ؽ=��N����z���M�/�ԺT(.p��l�ʎ���u�T;y����.w�����E��U����J|��*�n�`�����*\ӚP���C3�4��bٌ��%w.V�����F�y*ҝ�ƴ~�&��u]���I�w.%w͙Jh����p�J'�pƓ�Y/zu$5^���ҋ�������M��e?��$A������zDF�Y� єr$�w!��ԚȂ''�&NdM\Iމ�-
9Hs����wo�L[;x���{��[5R�E?	}/=�F��������|�*c�|�s���И�1������#�K�j"8wv+wnڱuۘl���4��MS'�2֡I��~�Ch}�f��OAyM����ciS��D�J��Y�	Xo�g��׌b5���8&�}������0mZ�;Ʊ��{�$��,R1�A\M�y�\J�����%dl���׃f� ���a��{�,�[̐Er��`��H�l1���{3�`��I�i�w^�3���ė�;��y=�jW��eL��󍩨lLY�k�]��Eh��[KR�˷��{��[+B�˷��o�1./W/g�y
�֬;��:+.^�u暷����4暷��k>�)0A.�fӘ)�@��HXw^�*M�CL�m|o��s��Ek�εu�˪w[�r���M"�r!�u�8Ʋ��z3��1!�C�*m0�ƾ�l��gg]����ן�u���],(��gumMemҹ::?��^̃���g�&]Ҕ�D�uV�!]ބh�k}74���qw��»�K�u���Y��;b��뎸ꆚ��0��/.${W%}1u[��l\���g]�.���Cr�IUc���c�t�8�a,�Hȵu���Y�oܽK��W�)�@&i޴U*���Lj�/���s.߰u�zQ��|r�u����<k�C[��MK˹|��u1�ގ)d\V�ؚ6�7���86v��۸;�r���g���Ǻ|}Ʊ._�q���C_���o��R�U�󔩇.iL]�XE[��(ۗ�Vp����\�ai9�oXZ����s��{g]���Y�����(����#&�:�ѱm�-b2՞��m�w����=V4�C���X�u)(m�K]T���٭�u���mr��8��@�E�R$�ܘ"�*c�\W�uw���w/]��Ĵ)��SHߗ�i�7E�m�*��Wwg]����X����)i2mW��Yڲ�(���ι\x����.l�[�Җ2�|��{5��aR�_���7ȳ.?�������é{���x�ݟw"�������^o?�
d�Cb��l~�F  ���(����l�nF  �&��f�a�y+�d�%�Ȟw=A&g�qff�	f�QH��5(N0�M0�B��Z'��&�G!�s!1�̆����#�̊Ӌ�-��̎���-��_a`	��`�p�7. ��q��(${.cq��q��(${.{q��q��(${.����_��	f�̎;�����e�'L�av��̎{�G!%N����0;�BJ�`v��8��8
)q��qR�[TA!%N�e�=غ

)q�����'��̎�G!�?E=#�}�I�$N0;�BJ�`v��8��8
)q��qR���(${�0;�BJ�`v��8��qR>p�	f�#,G!��a�`v<��8
)����f�QH��i'�/`v�����q���f�H��L�g�J qꊸ�Q�@���qO�D1}�+�am;�}��^��=7%#���{p �Ѿ��Ǉb��(��ԡ�I��o �fT�OD{�}h���l��6��}r���]!��ҧ�m+�`���J9��y�K]�\⬺"��A0��pF5�T�����3�\3/uE6�IX��,��ߦb�XuE�CD`9,w0;�@��RWDc�k/�Q��QW�>l��`v�R�̎�
�O�h܁������my�'m�Q�=����u.K*�k��*r��Å��WZ�:��%0=�#���\	hp%��4=��
��WR�jOӓ��@�jp%��4=��
��WR�jOӳ��@�jp%��4=T�
��WR�jO�ö�@�jp%��4=E�
��WR��?t��K�-���8:�Uʺ��.�y?JG�:��
[�a;?[��q���N�����+��.e5���aK�lB�I¦'��d���-�A'#�LL�-����:����Tؒۼ�#[��L�-��u :�]�t �V'-[d+���˜N^�t�����e*lI�m�/ё�Ҏ�Җ�N^�t6ŜN^�t��z��쌩�%��nIG�:�c*lI�m��ґ�N^�t��:2���e*lI�m��SYct:y�[4,R�:y����T��2[��N^�u�2���6�oӑ�N^�t��>t:����Tؒ��OOG�JՊJ�:y���˼N^�t����:����Tؒ�ܧQG�:y�
[�a��M��V'/SaK:ls�L���e*lI�m���#[�*F���6�1U�m���Tؒ�܏UG�:y�
[�a��ʪ����l�-)[��,��e*lI�m��#[�/ɔ>%Ө����ud�����%��ﲎlu�2���6��֑�N^�t��>�:����Tؒ���[G�:y�
[�a�����6��e*lI�m#[��L�-��}�ud�����%��߽�lu�2���6��ב�N^�t���td���C�͇N^u򲨓���%��<���e*lI�m>�BG�:y�
[�a���Б�N^�t��sFTd[��e*lI�m>/EG�I�-��羨�:y�
[:̖{~�1��Q9z�="��G�u>�r=8�������_���{�r;$�諎8��q(W��{�r�uR������Q*v@���ޫ�Q�r��z��*��-�\���"W��{�G�U���ޫ���T�zpm�{���}��z���qT�\�\r��z����@ɪ�=�{�}���l�6���ӑ���Wo�E�V'�Ra��{�\-�I���^e�ͨ#[�L���ޫ�3&ud�����=�{�}V���N&v����H��$cG����Ց�N>�����:��ޫ7�"e����f�>�UG�:y��n�7�"wt�2��{�� ���N^���x��`��U���ˎv3�)[��L���ޫ7�"e�����=�{�X�z�
��W�g_�ķG�����֑�N^v����H���ˎ�^e�E�#[��L���ޫ�3�ul�N^v�������{��Ǉ��ǧ4��
[yc�.��'����b��QVmS4'�L� 
AP�g�q��e;�!OT@PJ�\�g.�8��u ��h/�ggK`<&`
���Qa*!6�*��2dV�Y���u-�9k�h�N���Ő�+���/Z<����)��f]�D\b`0Z��ZLc�k/�[��mqo�Pt�	�iM(�`�E\C�lF��d���o
APܮ��x�\��%^�H$��r�K���Z�RAP������$���5�,��	���10Ş˭|�d��S��ԶL��������XmM
�P�V�w��]~$�R�ه��e�q��d��}��B�7��P�Җ�H�\B񍩨lLY�k�][Nj�@a�Fj�@�7�Fd�@a�F\�@)�P(��]aF*zƚLC)�����o�s���
�붏u5Zg�S�LC՘6]��l뺾����Pv�4�X��mL��Մ.xӄ�7M��V�P��վ�P0\v�QS��K2��	�w�4�hMٹ��}Y���h�Bٵ,��Z�1�Uԛ���	��<j�q6�M�$|��˅��+ʮ\X(�r)�XPL��}th�h��w���q�����,�]�P��l�4��:π!�4!���Z�Mi#1��e��Pv�e׫�Pv�Z�5�Ua|��tHޠJ�f�,Cٸ���e����3Lz�4>� �3���u�>�>�.�;_��h�0�)�V�m�ѥI�_�.�}����(F�>y�:[�t}6�+���#�pPv���{;��epY�bk�4��oǱ�Ø^�>
���f���i��f���i�n��BُT�¥�6���X]R��6���vuQ���O���8(�>����8(�>����/,�]}a���K_�u�Ue��b�o[c��|���r��B�՗X��Ec\��#ץ��.��uQyg�e��M���>����a�՜SrQ�b���-\X(�\JW�d�I�leB_v������)�,S�S�sa����0V��F��d�B�D�v���-+o�#f�`��ڗ@ua[ߚ�"�i�)~�24CJ��b��'b��~�?�aNO�OO��p�ݟ�¶�Cӷ�c�mt��}>?=6^�;
D( {~V#�=k�Ȟ��Ȟ= �Ȟ�)�Ȟ=3�Ȟ�<�Ȟ7� �@@��9a��m���8���3�($�������3�($��Ӊ���3�($�\Y����3�($�\����f�QH���	�p�w0;�B��E�N0;�`v�d��!1�`v���8
�>jb8�츃�q�}.!Ť�0;�av��8��8
)q�-��츇�qR���(��	f�QH�̎��'�G!%N0;�B�� ��(��	f�QH�0y'�0;�Bʇ��8��x��qR>,�	f�̎�����0N0;`v���m���x��qR>|�	f�#̎���a�0N��M��&̎G�G!�C)a�`v<��8
)����̎���{0N0;^��8�{��SW�me�b��q���L�Y(F��{��Ѿ��҄b��,����J��@(F���{��Ѿ��F��0��Bb��?�q�n���}���x��XuE��`�`�Ī+b& �3�($V]�y=,���q����,�	���8��ݜ�	f�QH��"v3h'�G!���͇a�`v�Ī+b7�]Fz�6��mִ/��/ �T��
��U�:;�"�����ϴG����T�����hT�\5��
W;?��
��WR�j�gڣQ�r��J*\��L{4*P�\I����i�F�U�+�p��3�Ѩ@�jp%�v~�=(W����.�h�Ef:)�
[�p�=)[��K'h�E�V'�RakN���"e��~���'��a���I�T�څ��H��a*l��pX�luR1�v�D{8,R�:�
[�p�=)[��L��]8����NZ���.�h�E�,��e*l��pX�lu�2�v�D{8,R�J[b:y��D{8,R�:y�
[�p�=)[��L��]8����N^���.�h�E�V'/SakN���"e������'��a�����T�څ��H���e*ls�3��$��L�-����td�����%����lu�2���6��ӑ�R��R��N^�u�2�����%�����lu�2���6�iԑ�N^�t��~�:����Tؒ��7SG�:y�
[�a����V'/SaK:lsS���L�-���Xud�����%�����lu�2���6��Ց�N^�t��>�:�U��L�S2��,��eA'/SaK:ls�e���e*lI�m��#[��L�-��}�ud�����%�����lu�2���6�%W�m���Tؒ��_]G�:y�
[�a�����V'/SaK:ls�{���e*lI�m�ۯ#[��L�-�����V�ˇR���,��eQ'/SaK:l�y:����Tؒ�|���lu�2���6�ϡ#[��L�-��猨ȶ���Tؒ�|^��lu�2���6���#[��L�-f�=����0��{�G���;�
���ýW���U�1��^=�
�����@�jp=�{�{���\�up��R���ýW�����p�U�[*r=���=�KE�\�^=�
���ýW�睩�����H5�jp=�{�8*P�\�^e�=���d\*l��^e���#[��K)��ɻ�v3�)[��K���ޫ7�"e��~��=�{�X�luR0��{�� ���N���x��`���I�T��z,R�:�
��Wo�E�V'%Sa{����H��e*l��^��������=�{�X�lu�2��{�� ���Җ�N^v����H���e*l��^�)[��L���ޫ7�"e�����=�{�X�lu�2��{�� ���N^���x��`�����T��z,R�:y�m��Ï��Oix[��Ɩ]4�O�U���6���ڦhN�BA�� A���RBP*J��:��b��0�K�%�F�	��a�(1a��a�؁l0F�F�F�F�F�F�F�F�=F�����EW���ք����P��5�f􌨆���?�8(�󉃲?�8(�����?�8(�s���?�8(�3��u ��h/#�a�`��հ`0��T�>�c2r}�)�hj��CK}G�8��Ɗ�����m+߻��.?�s)��Cc�2�8�c���>
#jW��e�	�7���1eM��.tel9�)Å1PA�1P!�1Pv�8����+�HEo�X�i(E��~�Mt�t����K�Ǻ�3�H��jL�.Ox�u]����\X(�\�v,B�6&�jB�iBߛ�Nf��u�G���B�pٝGM�CL/���&�9�Ģ5e�ں�e�;Ƣe��8(�'ڵc,��7��B=�y��l웾I��ۗeW.,�]��Pv�Rt���.;���6�T�&G]G��ѷg6�P�=l��l�4��:π!�4!���Z�Mi#c6�P0\v�e��Pv�e׫U�PS_�w�M����n�n�2�����qPv�Qo�!9ä�1M��c
2�q0�XP�nP[7�sa��s�Ҽ�Uk�&�	C��m��v]��m�%#:d�����<E1�n��#��2��yH^ql}9>���˥.���1,��Z[Ӧ���};��������P0\v�4ewN�Pv�4ewN�Pv#U�~��.�p�q>��z��յ�U������d|,�}�A���}�A���]}a���eW_���C�*ӏ4�k��x�[��K<U�c�ʮ�Ċ�~(����.E�w)կ����8ˈ�X(�\l���8��f�E�S��ܘ��*c��n���B��R��'`M�e+��3m]���MYd���j�e�O��\7?&��$�+���mYy[W�0�e׾���֤�L�O�K5��aR�T���?����>���N�Ç������w��x����çӏ�n�O�?�������V�� Iݿ�_�33e��Z�ܙ�#��X�3s�DR!!���3�*<֤�[n��I�,yϴvg梹d�Irg��������o�7�q�7Rp��9\ycL�"��Z�3s��՝�ǡ�ۇ���%�;	�>�7 �L�*���5�t���܀zI�ԔX�%��ť��0kЬ��[0��m����)q̄os��"f�0�ٟ�̶�.���H�L��ޭ��2QY���n�KQO�H%ߟ����MՌ��[���U>��������ɭ�N�ZQ����QV�)T���W��ԫ��:�4n�L����SD�=���쩒>|
;E)紵����q�$��V�n�G�Dj(J����$T�r�J1ߚK�Mn��c��r(��ǋq��dj �u�m..������oi���s���2:��ո(K�M�t�P �.�ݝD(�b���@G��g�u t�U�����:e�-��}�/�t��M�i�<��B:�+S����hn�-~%R�;�L֒���XB�2me����ҍ�ᇇ��S�_*��m"������߬�f��[���% ���$�6r�:��W��6rª�MoQ|#' ��Y �S+�PԮ��|�oQ�#�7oU�#'(�aIJV곲���+��)��u�'P��y�ʧ �TQe�[T!�Y[5��bD�$�ֽ�^�f�6��@)� �"@P�0L:I�����O�����@���:�[��	��� �e{ 
��= i����@AZҷ���_�`��]�����Ӫ�İB�IB�#q�$���hr� �Q�$D�J+q%%�����o���k*��R�^e��4��R�lߤfs#NyC�>�x���۔�B8�+c!�@X ��u�����=��g+t�3d����1� �� "
5�V���o=�!��[�AX�D$�e=�۳ IQ����Bx+x=<F��e�Y����.b���ƀj�!���#x���;���.�������S�4�}�����L���p������O����&�$+�C�s�I!1�=7��C�sc`!1�=7�C�scb!1�=76�C�scd!1�=��%d!���sÄ,����1��BXO���OP9�}>:M�`C	`D����6)�%�!�c��Cq�< ��|�������� ��|J��Z�ť���S�iy�`|ϧOh��upi!bYD0��`����\d)�-v [,ǰ�'3Ky l��b9�}>zb���`�݂-�BZ [���2Z`������.-�-� [,�H<K [��X��x l�#� �b9F���r���� �H< �r�?ҕ/��k �3�1�_�N���w#���� �U�q��w&�g����(�_9F�0�r��`|�����1��c�S_9F�0�r����1���c$�`V��x �� �4�#� �S9F���r��`O��T �#wz� ��`O71��5�ۅ �Z91�v!�LP�b�91Y�!�A&�¯�ז4�����b�L��B�]&�d!��.���Yl�+��Y3e][��8�����{�V�"L/��n�py �� �Z�qm��_�:�\[E�W�� ����b݊sȵB~�1��_�S&,���f�	���o���?s��XjNF~��E����*AXe��ە&�jf����f�	��l��?|��G�G^jY&�"?B��k{�bg�ҏ� Q�f�
�����V�������B�X� ��B�F�:��-Q&��x�K!!ެ�lO�uKw�b�'�߬W��������������#0?{�`�y������N[� � ���#0?{�`�E�����Ϟ
��
�����ϞJ��J������N�fG�A��G`~v�f������t<��O�	�0o��eOJ�Y	�a��A������E�l5d�I�����0�����% �w$\n��R	�S�i�a�H�9̜�T�,��i�!��-T�ѩ�!��;�A12D�3`��`d8K�ͣ��@h´@X�&��q:�3$4�\��!:�3$4�\���!|��݂�qz�š�0CB3̵!h�w]�	��;F��0CB3��k�bd�N[��:����������&?2|�H�Y���T(�b#��!4�yxye:���,̐�s�'��Y�!��NUh��0CB3�]��2�׍���Y�Gg1�ŀ�a�n��!:�3$4�ܙ-CtfHh���Z��,̐�sG<��i�!��n~h����	�0w"�0��0CB3�]�2D�)`��f�;@n��\����cD�N[�s�J�Z��0CB3̝7�2����e�捄���tfHh���)Z��,̐�s{V��Y�!��ֲh��0CB3�mq�2Dg1`��f�[��e�Y�!��v�h��0CB3̭��2D�-`��f��@�e�N[�	�0��F�����an���!�k}����<%���S�	�0�=G�����anَ�!:O3$4��n-Ct�fHh��U>X�:O3$4���-ý�]V(tڢK8`��cEߠ]�c�V�0 �=�ag�k�������qO����q<�tg�m��%~Q��L���;���Px�:ǃ�.{i�8D~X~:r7ˏ���=*e{v{�i��=а�8D�X~rO�ˏ���=�,?,���A��w�a!����؋
�#���a\�59'{��8D�3~�"M�t��3�"P0�#�٧<�e��e�!��!��v�7 bd��[����2ոV�>�-Rt.��x F-���/dT��!:�3<Ұ�}��vX�j謆߿�@�Hщ�; ��9�ѹͼ;�D-�K��f����"E�7��7 bd�ex�!��@�8:�3<ҿ�}�!Z����H�B���h��b��1褆��@��Y����7 bd��b���/�p)�k%$�s=�"E'5�f�	���t7dQ�):����pIK�Z]�xU�H�9�w���D'5`�K�'ZT��1"E�8{��O��~������)]�V����eM�rU�q�M�(��)����;x������N?x����U���������m� ������k+y��Iվ�͎�>��bՖ�6��rJ$B�^H���g���~`��vɔ����G���dR9;ǫ%x4�!+�����uܓo��KL���t'�t'җ��p�	���'D�<���u�e�{뇢�LpMkBQS�h(���e3��|Fڵ�7��vͨs���Ѯ��|:�F0�-�ù~!�Z�8p՚�����I��*�V@�Rԭ������/c�-��r.�W"���Y��,�߳f�Yx�g�wWC��a�)�^GS�v0mZ�;Ʊ^2�+���`Wԟڶ򽫌���:��>4�/C�c=&��/�[��,�v�y�P�Җ�(�Mp�1��)krMz�]��<�q�f�¸~3g\��o�"��73������r�z
��EW���ބ�&�P�Obi���\閴s�����sef�}���:C��d)�ƴ	'��u}�S3,�[1<,�v+v�i�"�mc�&t��&��i�d��X�z�%v+˂[`�A��6fVS�ӻ4���z�9�Ģ5e�ں�eջ�:����u����ecY�@�\ߘ�!ͬ6gc��MB�����x~���Ϻ~���.�g�&�������8�vx�{��7���tMS����Y�t}������Д6���Y�K�!���g]��X�ox��j���.����z���mY��qٷlɟu���{�ɕ%��I���)J���cAE�����Ϻ~��]�)�jM�2aH�������KӪ��7�Ϲ~��e�E1�n��E�y��+�$Nnjl}��/������{;�PbpYbk���M߷���aL�q�����ߘ��7�����Ǻ~c���߈Y�oE�}�R\T�����.�N]�XE[��(ۗ�Jr����\�e9�o�_��[��s���g]���Y�o���(����#&��%Kڶ�1YpOU�6�?����+��h��s*���ޥ��.*Oc��f���~��6��~�d5�"�O)�qnL�t��J^�ܼ?�������i�Z�2�ʄ��L[��):oSbU�ؾں?��-��jp�h���Fh�ۮ�'�e�m]Qp��s����?P]�ַ&�:e��>��j C�0���)��Ϻ������^��?==�৻��t�Y����w9'̉\Ϋs��3ؼd�W��:U^\�ˑ�L�>��c+��w�>��;�+�6.�����y��|r�y���w^�;��yޣ=o��K\��G�����g�R�~�'g���=��%��8�&�O���X3g��NM5_�H}�ϗ.�䌋r���w��N�_A�FzquGN>p}#��~W����N���C��gq���#p����xuǏ]�7��M��u�d�??���S���c~��J_���eRɪ���a�;Jv}�d�D2k5�=cI���A�ʃ0ך%rs2ABFRS,��k����%����)$d$�Fd�2̍LII��L%!#yMK���"#o�y;ؼY�.Y�yX�y��9�k�>M�>4�=��.���_s�N(���y��?n[`�E2�/��3
�9c9S��s�QH�5an�e;'[�����������dKY����ɮ9f除
nN���!Q�B��֒nٔ��zNg-R�V��ʙ�t��mnћ�zNg-���̉���tH�?��܉�������8��
��}b@~�Q)e$�Q��U���,N��hI�j��Hx����ˌ��B�N�h^����{��т�{��}����ך2��;1�_u=�o�d�,s�7��?�׸�7����b-�e
��"~>ͯzn�z��Z0׾&+���[���Jԍ&db���P؍Zd��oʜ᪃a���mA����]��b+v{X]bb��8���EZ�I[ʓC��I�~����f�&�2U�v��3���>�v�s��T��̆��"DX�6ؽ�e��C��1�I����Nq�\H9����
����҂��O�M;|�v����ix��lY'���O4�ɽ���?��������S��_~�󟊗���O��O�����j�S��S=��.Ҡ�8�8��<h.�����Dh.����2��Lh.���R��Th.����rq���\�]�?��<��?��<��?�����e�.rqs���\�\.�"7��������.rqs���\�\.��~��"3?���2��2������E.~.�����_���r����\�E.~.�p�K��%\��r	���\�E.a.��Ų��.r	s���\�\.�"�0�K��%��.r	s�ċ\�\.�"�8�K��%�K��͇�W�����������XK%�?�ӿ>~N��Ս��O&�Ż��N���.׃�޵�"=�L�e0��D�}�Eѕ�v���;����iH�=���s}���U o�`S�P�����6v�ھ�l����kU�N��k�taF=�#5dB�ţ�ƛ�+S��齫|L�{{y�"圦�w��y���W(��xEɔ�~^Sf��v��K�|�/9᧟7O�&�O����Ï�����\��Ï�?r\��������y�c�C�s����?����>߲ȓ����I4w��>��������wcV�������z�~������}~�8�w�=��H������>?�[^{�������I��B��O��~�w�|��},�+��I���/�}���L�`�`;�Xך���oһg[��㧧�c�r�c��������5�����߽�>//�T^�B
W�K����ֻk�/������ߗ����+�ɮ\@nrEy�!^�@_~(&P��ʭ�P�\�h�
�V�0I�X����i]䁎���;�u\XM��� 篅��q��症�	\XVTӗ��~aXV��˗u��?{=/?L����Yg.�>W���j��Â���0W�������?�?���s���߆�O�3���;��c{mkbҲ���zy���|��^�H��͘<C�.�h*M(��i���ug��CW�sc��fjl^|Ӷ��b�k�zN����~6re��r��X2�2lb�ֆ�<���+ޢ0���o��?�����7?6����?�4�^�/ȿ��V����x���z�P�[�d�:����L�gL�ʦ�}�a�N֗U]N"�����U��,�r.�����e5;��^�y\�������/5�A�w���a�Y��>���+��>��E!^�����W]����D򋞾�����i>�G�T����7PT)Ϊk�kh���ax�2J���?|���먯����7�c~y�Ο���/�U����8����.�������zA�g��>�������������7��e�"�����u��I�BR��U�,�O�[eU���CYե���|=kJ�C�%�m����416���ʮ�b3�5��Y�&󽎗������K4�闾�����6��2��?�����g�M�
nM]��)�L�Ug[t���|�"���F���_�RzUU�Pʞ�P���i�*Y����o�.��T�X_qNU����~�K��aF���ܾ.L��:o5�Q��T��Lj�)�2iE2���(E�,h!�����Y�sQ�}5S�5��Z����;uOIiII��2.ǺY��w�:X_����@��=O�c9Y
XQ������	?��_�瞚�:<��/��}x�G1%b�*��
Ž����'C�"�p�>��5E���lSu��������{?��%N�Fvf��:iy��$z�Yyƕ�]J8]YI��j�{�*g]^b�{�w�K�������we�%��Ub�<��w)4OI��ߕqy\�J�K�'=���wy!�G*����T]��L>Y��..)tU%g���]���J����v�u�/����J���/��ｭޅȅ˰s6�IE���Z���]|ֽw>�Jc^�&/9���yB*G���\�9��,�����5ϊBxy�zy���f���My���ֶ���f|����o~�����>��NH����W�)���"�pQ��f��}ms{�:6�T�s��t]E�؏�����1̎�QW�7q?�yʟ*m�V97���WU�%��vW�B�=%3�|�eQ�:��EYXͪ����M���o�%9���_�Z[�˂�K}Gt'�1�\��x2)_<�}�㻐�VM��Д};����Z�419e飩R P�f(S�<�N�1N|��;W�8/u,���rd�7�OA���%�,ޗ��^��=�� UV�9����?����{uQ��sH��(���H�}W��u~��'����{����#T�4�`SH�Rkb�LQ3�ȼ.f)7�� Ǧ�}NJD�f�=������/���W^�:��oR�~
۟o�7�.�Jn�h��ސ�9�����C}U���dR<�)&w�Ӑ�땆��ڮ��9q�RV�H����+�{S-ն,��x.��E�2�n�\�谂�0n�'/�0�ۮ���,NB��Z}��_�LcWt}4��sB���1O�JIp
&F?6�,6�4���c*&��R�`(��叵���e�G��ԫ#�c��X���������������������������?�=UU��HQK�%EY�R��|�K�19�@�j�/X߷��ti��R��KYP��0���K��4�������\_��>r��8��M7� ���_�C�/�P���|J�+O���I�y]��r.ɜ�z�m���V�54��F�\PU��X�atCr]������
�+�ϵ7��'y��j`Q��q�
ݵa˻6l"���e�9[��������"r��?�X�e(?M�P�����E�>Ԧ����ާ �L^��j說/�&�"N�h^�/g�¢��yH�8nZP�6��ֱ/[��ľ��[�@oqܜ�|���;k��s~x�<�!v�s��*M��������U"���/G�D��"����7ԇ�����"��Ţ"J���.�D�W�*W��.K���P����a���)|=3��b9M޺�/��Uӿ��'_���s9kL=���WQ�r�,H��C2x^�'���r�@T��͏M�~O�_�z��y�b���O����gT��K�u�L'�/�BN��H!c�2H�s�nRV}�j[�Ɨ�\���g۹��I8{�����z���\\,l����,F~e��o.�D��ϖ7����!/&��v.�Oϓ�\�翺�0���}g|����6��>�F��C7��qIqN��.k��x�p0Ա
���/	L2$�˃�,Q������|J>���+�>-]z�+*|$�չ���w��B<��]W�R�V�kr�sEi���4I|�]w]��vV
�:χcA�ݥ��4�����<|�x��$�;���w�&O��yx���w��6��?��~��*�w��/?���,���r������қ���C��/~�8<=�׿����镞g��~�����������ߎcV������.��ǧ_��������'�����&� �3�c�� �%���c�����O�n�~����~����`��_�~s^�����������h���3����" �0�z�,���Ͽ��sR�[��{������:��ֿ���������ۼUL_�˨��y�0�j��4������rU� ;�AXy��a�]��b�ee|]ξ0�<�S۾����M�窕�����=T.���_3G��q4u2��ǜ�>��+a�U��*�u��5-��
���k����Z���֩�)ƁX� 5�b��^wPYU�ɨ�������k^̓�M;�ܘ�u&�mI���Pn�$h��|���:���?�a�_�}V�z+� ����j(ݸ1U���r$b��e�����1�i�u�w�+K7xG͂�h�C9��C����t��뗗���+g��e����V��˃x�����`'T�/_J_�L7��Q_?ۼR��b�F-+�/~q�זb��:����{��!��K��+ҵ�,:�ɠ��?K�@�V���f�
���U���b��B��f��E�1�Hq�_w�ᖣ��*09	|O��5�>�&�����_"��_���ͻU`6��q�q�@�ծ���$%�GU`b�ש܎�X39|D��-p���Z�}�~���)��]��<>j�(�PV�]7�F�̣��^̹ ͋0n�t0�G�@�z����ō�8���_ǅ�eQ�8� ��[Bǰ7���S*�<��+N�RC@W[��qW��J����q����C�nPD�vʊxc*u;�ÊX�,E�����q�����qo�J�Wz����e|�ٕN��O`�YD��������+6`AU��^v��vG_�KC��:}mey�6�U���U�K栫Θn�糀���i��Aq�mÛ� ��;ZH��Wi��k����ϕ�;�2]�
��<�E�-Sq�r*�ڃ-Hx�wP{�����:�\oЊb\��5ӟ��'-[��`�%�Ek5	]��՚tS��䅮h��������1s� ��������Z5ؕG�U����VU�z�J���f�F};� F��ʁ�y_�U��e7��-��\w:�b*��֕��[W�z���t#�����[�������;���5���o�s}���/�?\'�x��Yݰ��,=3�em����lo� {��z�̾�\o��|�q}�.w��C��T:f��z�NQ��t���r=h9��t|P�M�.���Jw��t��|����������Y�(��^G팳7�Z�<��;� �کDW���譢+R����VL���EXŐ������):;G`��nrv���s=l����q+�t��;E/�,ZYntS�sS���rmV]�T��+x'�Yl�Z1�5+������dI&_ï��]����Z��9��A�����G~����?��wWd��@���;��� ���IG�0�j���tk���wq�#���"uG��
g��S�>-e[Q/{�r�O_���eڵ�W]�Vr�v�i|[�,Sd�4.�t{�}��(B]�BǕf�q�zM`.�p��Hj�,P?� �mV���\7g:;1fA?�ۭؽ�u'���n+ߝ-�+�7�4���[����.�*���7�M����oy����/oDN�Ϳ@��s���ᤫ���U`�������i��*�UR{��e%�
* OQ�b��tW�|�\����#��R���6�'E����vr-ܘ����n������̆o��8`V@^V�m���M��0�q_{�� wK�6�ML����R�T��������0Gq7��F�gk���mk)�1v��t�Bz(�Ps�(�}�U�J�U%���E�l��1DѶc-�NsW�0`�㚲Y�xC7�l���f��hsx�,��C�e.��0��Mpz�^���{9��)�8�-^�V8n0(ja�y�T)�����o>�����Q�Ba�#�5�3,xuvocE�}ٴ9��2�V>.wF���V� ׹��!����se޷v@�Lq3]�[KY�F�e$�\�ӛ��r�?^K$&��;��7�o�+l�@U��SuӅ�BL�@^���ʮk�%����Ç��y�7>�}�5��������c��s��g?��i��S������� PK   ��V�4!V��  �  /   images/1efc6cd5-4b9b-47ac-a031-8851919f3fa8.pngT�uT[]�Z�@���V���ݡ�-�ŵ��H�Bp(���=8w��C��o��G���g��ߞ�='�<&�/p>j>?_�@�}���/�X�����)/��b��ϋ�/?Ji{�]��c���C�d��Y�Ƴ�IA����N�&���^r�x�ղ���Ӏ���)��t^�&�ʋ�袖�>\hG%����,;�F*%W}��V�C
����ů������r��1���gi���A������Օ�Q�ϟJ���d���R����k�ג�sM�4$2����������ڸ���!|i6���� x�o@U��������:ٷ_��N=��'�y� =!����^��i� ���T����?{���$ndl|M��@}ۦ�|ŒYZkR�$9
�>|�\�tE��~��n���G��-�������L)�ͻwl� 0�G����է��5:��H1ׁ#�˿6:����8�q|}����e��r��}��Q���J\�����t��}���������j�cv�V��˞d���{��v����'\*��C���A��E�9Cf�ùh��5g�x8�Œ�Ds �����7��v����cK>�<B+��̷�k��"��!9*���K-�%�ԣ&fc��	��6��Pݭ�S�MI�z��������R����i1����,ק���zF���	V�WK*�b�l�j�2?�1ߟg�aT86,�h�8=t+�^hH	h����\��q�3������f���o�銧�S)N����J�B�U
����a�.�f!^��3��=:�����Ꞛz�:�:��H͎(A�Qe�XF����7�Gsq��u���?�o�
'/J=V��I�����H�ۧ�ȭge�4Q�"�	��Ѳw��Ld�ځچ@� ��SsЍ�I�a��rU�(��7��V�m86�p���4}$�Y����8{=����bǳU�N��aA+�-D�	�e���{]��~B��O��
��H�@�I���Mu���h9Y���NM��sqvv���X^V����nk��H��5���"��߲f��%w�-�sd��&�����b$��o�k��.��[��c�������Cc�F�'):���GP�1�ܝ���˨�޺�|����{;�,f��:<��K@[[)���+�O/u  S͐�5����?j����݋�.7���.�x_Qd$A����������j�-�0u����䕀?f�u�ً+YPU7U��H,?��!<Q��Wk
V��jU��e�����H�b@�p�;�Y��z��~������f��\%t:�C�h��}����a�$	��PS-�!�32<�}u��ʤ.�����Xv�x���A��-y��i����<�`���:��M�/l�6NƂ7�&��(���z/��V�����`p"j���G������iGd��H�#G	R���$<�����f)`��<��=Q��"�0��"Uz�`:Q`���G���r�N�����^�,��_�Rڎ���ʲ�_� �
.�/]S�7(�b��~kk-J���rU��xK�� ��g�����l"6�v�}L���s˼7��������^�Q��=s�ͦ���᱉��Q��y�VK� 4v��A<M��70ƫ�)V�Z�����o�N>݅��XO9�oZV�����~DMBJ�@�h\�{��I9��)�����k�2r�,E��R%'�Ԝ�&��	M.������nBZs�WO)�EW:�-��{�@�&
�c����乏1��c�s��j�8r`^��n�sT���_��]���6�x&�#>��s��F����NO���>��~7�j��d�Usڮ%���3#���a���C~(�"ˀbsq��0*��6-��hB�2��������R#���@k8M��O?�X�EZ�O�@螉%�U8�S�֜q��mY��S��u�~��PR��(��d�$�Ky��7��Ȥ���LA\���/���1y?�a�lJA:���z߲X�%C��|������l�A��˺-������:��ޝՖ��>|����m��?P�F�M�q�=����42�����ZGBU��J���E�c�<�~���3���Ws)hk���1(m��s;h�k>Z=�'�.�
VS��]b�UU�� ���/[��'�{����{�4�>�:`h�?9��_�U�p�.H�Fl���Y?�M�K�.X%]w����������;��	��?A��ɗ�k���4��3�� y������>������#��5ڳ1�Zqb4{Fڵ�C�s��z�u	��ߙ�����!&ǭ��y���Q��s���`>�4�g6��^�"�����\���E��]�u4D\�(,&�Ե�cl� o��o.�B��7����Ky���;ٳi7D�˵�/h����%����'*����J���,�^����}?[r��V�u��
�2>�=BU�iT���ʻC0��/t��4�_�8P������[���6T�������v��p�=ݒ�X��*�RE�U�ή����3m�,H[��Ê�>���KmHƍ��`��K�H`����wd��J�! �R�<D��J�,m	`��\�YоB�^�6�:�X�
z�c'p�����^�5��������(�3�]J�&��v�VQ���k&5dr<غ�/˳l�>n=�h�k���d+���%WYR�S^^���bL���)�C��2��v�����h�_m/��fH{!��Ǝ�]�0��O, j�� r]옂p��m�hI���Q���*�vq�E��H����)ƴS��N|��g8�+c�����-/8��x��6��0^|�f���~>��i+_櫹{]-
9Zˡy̽�p�:.�&v�=18�
���w�˟ �cb+�� ̝K��,{J��1J�T4L��`��p��E?aӧ�T�h�]^w?y�<�$eG.�]���Y�~�M������8&�T[�%�D��N�xr?>)�Ԓčqx�;�+:H�����o��HL�J{�g���,,}�+&]*'?���sr�� ���zzkx�U���Y��U�,���LIawfc�P��3��;?X×�1���<�O��]>�>���.�-b$�߮�;��K�ăKg�,�*�}U1���iu�da_X�l�n\p{wʸb�Z�_����=!�k��v�.܏�SA�Z���:�H�\��x�^���W���s�������y���fzK�R$��c�D�n�c�%��b����{�����r���sdb���W���?	C��S{����5�@�g��Y�(�����C��F`�.�%ےۄ�Ǟs�M0���|�r=�W����k��HC�n�TV;�f�3<q�H��}�1����CV�����]2���J���-.uU$��;(Lz��f�L^��ĔH�_N�%�o�/��OI+R����km��9턞^N	����**���o���6�h*��s�%x�V��h
��c��G��*�>�t�R(3�G���ن��k=_�1���_�:<ff�Q+A��l����:Lk�W��.:�%l�+�7���_$s���0.m�:��BB{��pO�a���0>�m�t1�C�(Muؿ�-�t/��2�Vbh�\�s��,ߝ�2r��"<�IC����F�."rc�M��,�<]��)Gl{M����-���$!� ej��-U�nߒl��J�#���WM(�K��X��d(�ry��]9[Q�Q��Ao�u��wI�8��ZS,��R#�{8�a����qEj��7%�|�J���� 
o\5]�ӌ�������.�@-3�P�P���
�mNn��P���t������±���|�'ۮ�C�#'=ɔ���5�.S���S�V�Ɔ1���������?��%�m^��z��^�<n� �*#�<���p�v���a��P�3��*�����1�X�����b�Z >.$:������Ǜb%C��V�!����n���-a�'ާf��X�K�b�A9Ec�3�Kx��Y9c�m��DEzN�X/:��
�\k��~�*�s�ú����dJf��	�8v��mY\�[[�s�|c��� ��o+ahBko�>�_@��d�l2wۡ���^�鶺`�^6��ڪ��4s�,�ᢟ4]Č8T�e
v�|�T�D���!q�6�ݗ[_��ϥ���ǐOg��v�bS���2OW&ә�i�a�##i���?_�:�,+/��	alP����M\�!:Յ��'Y­���.<ݢ�U`Ax!h�f���S������ާI�)@d������T �����21�
���
���|�%��n�R�\=�X8A����"��',
�ms|�r|l�i{z
���*��B�I;�$Ҡ�d�(�B9��L>�J�{��Q����1|��~��T��P��p޲��ۨU�ɉ&d����g�Vq�;z#�CK|&w���i�F�%���b�Sp��˘�SQ6Gfc�^��ζ�	ЏZ�;����x<y��_=<qi��^�ݗ.-� �л3����!���c�֪���܊'6.��p֙�2 =��&�'�B�)_"�Ha��y��y��6�ҥD�]_�7�x����%��ܬ��4"�\#)�2����Q�u^�����t1�'�1F��ᅯ3!ej�}�N���Fy�z�
���l����3o�A��|�pK�\돑vW_򽡳3����\��]�o�=|}J��E��+��a�o[����?'���F�oHZM^���0�qj��q'1Y��*�ƶRbIL|�5�z~UM�PC=d厑��g�~��4¹EB��YS/^ё_����c��w�ÜcH1Zz�R�ERԸB�����;{=���F���e��)��(���24���B$�mj_�K��-16mȜ�ʤ��L��L��? s�Xct3:�Dڼ�?��xS�}�`W�P�)�2?�w����`�_� ķ@jt�g��� Z�+�@LJ�s��3��'SsbY|s&���{��	�@��C��-����}|�B�죽�5����T���&��.;�|���^�Ƣ��Be�v���74>��ɇS�����T��� W�Xoy���l��պD��a�dg'C4:�XF3~��7�p�,���dSW�X����1e����h����ziP�;��Z�$�T�����K��N4�˪/K��"�]�N����x�԰��i9�cH���`��\����`�o17ޓ��$/Q��Y����B*��W7���{�U��,LN"�4f��r�� ���a��xël�b��Jp"ҙ�Y����H��T�Q(])�_�!���C��+���^���'�#�a������2��by�����Z9 L�hC&������ݹ3O�����d��q��=욅8k��P�	cGM���ER_ހ��~b���G�K����ۺ�;Ղ���Y�Y�+�{�@�S�������-��� s_m�{%��T���غ^i�3��?�:���Z���9H$�U0�<>ݽ��U2�K����Ɩ�7�K����-�jo%�3��	j>����	�8R�[^����z�Jt�Tr��.p�lo�<��z���J�Nڱ�m-~�Sh�[����y�3�V.�F�a�$�\�!����"���=U���墈�O#���Ѧ�C��fgg��hK9�f���K�bH�X)�� �� ��2a��D��.��?���Z+qJ\ԟg��[�nzpD���%�� ���X�М�[6̦@�GU��P��HL�e�z��C"�!�v����ю��/KBV#�Ds�[�z�Qw�>T��伤�#(yS��.�Si�^A	E�s�>�ښ����ϫ6^�t�������.������8ZRd]�/�]��GW�\�"�C�=>��ل�!�O�*D\��f4���f��ɪ��|��FB&!�[���,Gd�C
P�/�=E'�#	�~#�,�����^��q�,�DU-��24Io�{vX
�־��b3�]��2�Uc��G�t��>M���glj����9�]b��X�to$E��9U�O��Z�B B���B���Dٖv%ܸ�����V����c{H'�*A(Rʀ��_� �����Y,�(��ˍ!�^��0�[�k�eX���M�7�9�d��B?��\w����J^�G��0�TWw��[m�yS�
3M��/k�;
V�
�w+���O�����-�m�٬�~EY��Vmʛ�	�-�]���$"xc�k�&���.��Wυmo]]Ku��j~�3�=v8:A�4x;�1le�>QZ���;>\�;�RA�cr��ڢ�=;T�d��wR	,��U&����{�lX�$5�:m�ssy*�p�I�?��Ĥ�J��jx8~�9�L�	����p<$�hU��H���[��d�[��\��,�s�M�ԴI:P�t���T�#i,1h"��2�(�����D��DH���ͣ���^+���,D4gP�1�:0|և�<�|�X��҉�6A7�8A�ٰ���>�8:�6���*A��3kN��2�\�J��M�
���r4�7�-��4�7���o,T��Ҧ>8�y�%ld=�
y���II�٭�AX��?����߉�(}{ч�M���I�?�=���!�W4�F��q9^��̭�\8�@Ӟ(� *�'@b��d�y�^��h~��'���^zC�G�qye6����`pɵ��M��<��>y.���x�+:��� A��Id�<�� |B�~�/�%���]+��K���=� �;9K�� -�)��!20n�h�������}�t��D�?�镍��v���H��l?/�N����;bI���N"�bq��V~$F�4������Ч�M�f�Sf^���@-���U�@�8� ��N�j���+i|�T��/�R��Ĭ�j���wМd���2�O�ڤ���{�����8�E��{�V�1k#i� z��Oʷ�
������l;V�:64��E.R��r@�g�q���chK�C�m��J�1k!��ӏ[��ӱt�c���+��0X������H�t����W '��3��-Ba���ƈ���bk��b�^MÂf���JL+".�4�7���_:(���?��@����$o@�-�a��>Ix0uT�йȄ�5�.4��T���u��l�n� ���h�|�|�6&h��#�JQԈx;ʳ�+������D �gN�G%�Hs_5�12����SX%���A����}���GE]x�N����+�E5(x}�� D���J��G��C�i t]��WD)�{��%�gə}ud�޵h)��Z�u4���5�6���@�:-eB���?o���7���-~v�Mr��tE�k��qŤC��Db���!�z�?��bA��o�gx�C�== Cឹ�מ�Jg�����������*�X	��d�tK��x���\��ҵ���jg�|�����W���|pS8=��t�h�լ���2e^bE�Q�7��PH\��E��*��x�&_Y�vt6uY�g�g}ޔ�ȡ	e%�M2x�������9��HP���������Mf�,9��1�#�3�(k����>��LK퇣���/��3j�Iuˇ�O���%����c���<>4ޔ��w���)��<v]Y$#Y^��ʂ�İ-
�ݕg�+7.�]`>E�%mYU9+h��2�s���:i�ڦ����K����ZV�>�ABc1��?H�޶������޴~8pR��#7���~�Cu⪘�]T/��z;Q�n���t�fq�[Vv4;0]����uk52 ��6���`f���@��^�9�nA��.PhM��F��r�P�>��8�{�:�q��8qS�Pz�����(�X�կpC�olң��9?�&��>����C"+&'����[��wM*߬=���ͷ�^c�iH�����ׯ�9Ȧ˵��9������any+�{�s�3��8 3Ym���/|$֫33xf����+GK�Cojap�M�������o�3�E:�w �����~R���+`���k&�K�o�����h$�f|YU�H��N���u��?�xg���EH}:���ȿ>� �"$?��_-�AP�U�ŻdϞI���s�⽼v�n�sy���6�C��# ��"�K`���d�49�c�{yd�Gs`p�4�~R����n�����7k�"ݑW�dc�AmLĪH��)����{��G�8Y���}��&����!�P�x�gNce�U,u���T0���sj6���T���0�_ʚ��ﭻz�p��%V�3Hg�����0	ٕ1o�W�K�;�ڑ}�e0fKy��,J>���-ב��3���1"�?�v=>*�m��ěMr��2��V��?�`.\���E��1%�����Z*�EJte�*��w��;o���?�K����M�X�#h2�[Ŧ�՚�;�&*.p7s�(ɗe��.^ XKc�?�<B���8㰠���q�:Q
�@)吉�Z�M����)��ZqAl)��r���b`�q�O;2���l��1h��|W֌�Y��=��"�0Mem���gL"�T��l)��0�a%�������O����O�1�{�$�*)�
��L$����|�G� 6����$�w9��qB߶ο�_�7}���,��Ru�O}Ȃ.s��M��}6���Ç`�s�H(A���s�,�a\oUؼ8�w�Zs}G�DvO&�E�^��`�Z��z�'$z��R�;z�5�]��"�p4!E6��ą������m/���lv���#3lnnS��`u�a��U��j3�8*f��KcfUS7�ܑ�̗0�64��bcYX�>g��a:����Y1�Rd_�-�C�-,�>��I�T��?�~3���k��!�Ӣ��a��R��`$\�	Pk����-/�f��Y#�&w����E�,������G����������� /�d�I�b8Z�sz�Б���L�����v�|��ڱ��z�����{�(_q�+�/��:h��H��j��'���*��������/UE��n7���KpaJ�4@D�%��Rt,����u'�Edo���xx+��rL�/�lHX�i<}���t ܿ~j0�[��a]�g��8�%���_�M� ��X��ua��I��{�w<>}	vb,v�^����30I#Nw��^���>�C|2f���[��H'D$��N�Ǽ�J��.4���^m�7�]����O�/�1#����bw��oW1��D�3�_���ZNI�>��V��a�_���K���6��pk�♤Iha=��U�$��^-������[��Zn�mb��k�"�riBe�A��?���>��wg6�:��Q5�@��֋���<T��N��d����r�S�� �7��J�@���r�V��0'�o�H�� �@�i?J*8cVe��?�K�q��{GO�t�L}t�&���$zq%��ύxݍ��!ak�Ӑ��D$b��c�⇊�����!q�����e(�jX�雱+���LGĿ��36v\��NU..SC}sX';ܴ~օ�ٲ�V�Q������]�6(mMV�E +��dtŶGʢ-֝-�U�p�o xO3�<��JAyFu7NDI��2����Ü��݌f����+�vuc���#�r��G�r8.|�>_���Ȯ�P?jh�)���е�})"<ԁx���&�}���-9�����p��u8�%��Ra}�䋀���Rk�'Z�ׯ�������oz�(i��WL}u������tW/φ����5BtK^h��i����~�(l͑��3G���7K�j�ꭰ�:7nԴ�ݾY��O��Z�������V�@�/��b!�L�ĪZFHLuQ����B���O��;�ҿ�7XS��W8�6 ��:!����Z8S�6�Z����d�		�ই��w��Si7:��b8
x��o@Kh�z��O�v')�9�����P{c��ί��B:�̶��]밢�Qj:=�KH�r�>Z�����fAq��+Ŧ":���ψӵ?>�{�M�x/����Egb�)m	|�߀ʞc [y��ߋ`B�M�Z«�Na���g�5/��	�Vt���"�R�x_�u�skn�9]����ʦm��R����.�B���PcRh���_/�!�Y��ϫ�����3���ƀy�xQ��VR��E韱1�5P�R���Ҭ��I3�G�^Ď�MI�y��!ȧa���8+�����P�ڝ.c�@K�b�#�c^(���n��=��UX�_�b=�q��U(���
E&(7�˛�ٕj�S�_���p���4��o�^I7�P?8���#��?��x�����i��q+z�+Tt���@�V�R].'��]�'��ب`V��B�#�j+#��*�1�D��N��XN]��~*�J!�E��ea����'>ǣ��n��� ŧHC����׺y9�"����`��*��?=����j��N�(Y�n�������K5��������C�<��{��E9�ȎmR|~G]�m����.
�˳g��,6�x��R�Iv�t�ժ�3H��Lu\�}��;5�q������$����SӾ�$x�zYfo;�fo�1�F]�,�^���� �d��\*�2��-�~��d`= ]�=�a��!"9��Q:��9�7/��v��8�N~2��J1��~`����9�}�"�;�\�H�4�`�R�	�v_�qx}�w�Sڕ��غ�V~{sy���Sp��"+����썸�z�*�ou�-i��z��?}�6����/Q
<w�Pc�W��Q挆ʖLر�����m[/��"�/��VQ�No���@$�\�o�x�V�������,�����jѲ��!Eu����_m���#�%­�$ZG���[�&4�2�'�g��K�k�6س�fzpڟ�~�!�X4�I�hKV5��m�A�aW!�<�pI"Lw�M!U�Xh�dfswl�l�hlv�24���q�ś-�{~Q�Y֢S�䊦l��F�����ѻ��ɨ;h��#�(��v2NG������P����@S�l{��7�n�rezu�u�m �z2�a��$0�!���o��fl�,�?A\CI�{�~I\:rZ9��1�HkW7�	Q[��u�V�
��4n��|��#�Z݉�e�v���3 ��t�_�94c�O	���0�Z�`�i��x�/K~L鑻;��S u���yS��q�X��L����p�<��_[���dq�^`r����|ڰ0��|�]�c��ފ:ч�޺eܰ�f~ǃq?S�+7OO�6�D��{�\�w�\M���B?��p���_@j�=NBL�pa#V9�Ǜ�(�~�0�G�r\O�P� y_�����q[�c�;S�+�[6?U�4�}��T�7�O��%�Ȩm<i�l���9��O{<N�ó��<��[�*�ѩ}�V>�C(Q���6-���@���m$pL�L2#��[v��$�!8h���A�IP}	/��X�F�$b��b����$&�]K>��5��߬�%������<����ps�İ��y:* ��W�C�D�K��g(�Y<初J����15�����}P*�6't$,�R��ҥN~YM�f�/��m	M�.�1K��Sd�uRy��K:�]U|Ug��%��m��.���R"�ƒR�ŏ�2f��;�j>�`љA��
�r��?�f�O�1��\]�ʯ]q;���%�����ZE�D��v�*PY[����꫉6?N�4����dt�V�K���3�C���[��^u�/+�y�0l,3Sɣe��_"�l�&^�\��$7ԄumM�Z�(a|����x�s]*�D�;J��u��>JRD�&[j�&u?�Oq�tW���[����%��e�J�7��oh��I����;�b��lk�}��9�RΫ�PtM�����D�޽\�m7��JV��Ӻ(���#��8 ���KkGb��Q���Tا ]�|8	Ɉ��QLL}AP!�2?[�ዕA�dHB�'�"Ϛ�.#�VKD�hŧ�������̖���qÍ�_S�^�"��	
r��~U�4�� �\0�r�6!�*�G�I+��~1ub?�OG�;�K�I���^{o�p ��9Ֆ>,�~X�Ǔ��~��/d3�lI�*�vT�	�/GC�,3��Vq�m�
o��)AN���/Ϩ��zU�Ι{�Sny�Y�t��_�㞃'<k.aD�T�ҰI��Fҧ�A�/i���W�iRn,,8L_�h�j!�'W"��~������}�+V��?�L8���蹐W'���l	.����k�l�Yz�9���w))Plu%����ķ*
����\!�+���ɓ��˂_:?���f�؛���5)�R\`zЇ,�:����>��$�vDr_݊��M��mp��#�'�S)���ѣu�/_���D�1���,)��H��ԣ���#���+�)���H�P���X;7�V���w'!t�,u[�#�H��O|�^?/���@��p��E�d��g��D���|\��
�L<����* kT��˓Xa3M���l�/|Jؿ&x�)�_��2��|�Z���7�~��5$p��$�7���U�ԗJ0�l��~�t��K-�|�#2�ڙ�%n܃��@�]�:�Y��>V1��\�ۯ�&��׻�����_AIP���pa�7R��n#+'���xc�͠/ &b��~�6���8��(�7�/>$��3-�wR�� �/$�ς,H5O��|��A������7��D�y�[��cW����°�o��տܾȮ0��Z��[��z
4���c�8|��:�Y����O���sE �+6��H��[�����ȑiy�.��7Z&tuǴ�P�R�.��O�\_��d>��ҕD�U����:�}�@(��l���<��Pp�]��������>]�1NB����V���K�*܌o�El��c�W����w�SvT���R�P)���Ħ��YD�O�n�<5��:�"3���	��g}�%wy��4V%���|M��x"��"<ҊF�u5�����6)��Ӵ{�\�0w��[���ɯ��7M"�X7{W�a67|�E�ul�S�����N���D*��F�v	�W-�@e��#R�cO$L���tŸ���ޅ��(O�]٬�m�B�V;םP�^=���c�=�s�@��%�ESU*x�fv��r(�ʰ��]ywƘvh���xP|�n��9O�`�r��R���j"'�E}��bf���8l�'���e�gz8��Z��`�lq���q����;31�|����C�W2�2�����4WD�*�J�Ri��a�=G{�G=h�����>���m�"����[�lC8���dc��4Y���������O4�Tc�5�ԣ��%�~!�IePH�3�g��Λ ����*�Q'�E�����*p��/ʲO��M��uП��J��=�����1q;�Y♆tq�¦��Cg<t:�,e}�돉���
!o�V��|$n��P�H��ۦC�8$~w/�1Q�%o2�xk��.jl�ӿc�/��G�3�\L�2�Cɻ��ո *��Ɣ���*~�-�D���T���z��w,.�גLẑ�blUmV[��[�}�H�y��|��Ԯ��({#%+<���,���:��{���:U��0����l�GRF$�O'�}��L��׻���Vh��e�ukc�7��z4��O��zi����
Ϳ"�l!י�5�I"�����o�`��qa�������jz�D�kݣ����f�H��$v˓��g�[�_�}�dUr�����z���F��'��A�$�f����4G+	�,OF-f�;��F���F}Y�my�]K���n�L$K��MU�Km�ZW��HCS5����J��1`H|ُ�6��2�3w�d߄�e��B䜗��k�g�NF�Z ����
um�:*�{��+X�%�_j^�~��������n �O!�V�-���q���0��{�%����H�'d͉��aBEA�M%Q@ZӇӬJ�\ڤ���,+
������U�@W�^�(�~{�K����T@�h�f��q��U�B k�����fa�!�/E�V�'��Ia����S��oˢ��W婄��ݠ��{��`����6]��^�X0QV,�?�J��/�m�(ɰ�9v�d�4N.��'��nj�3�I�1��#�w��Nk�P�4���}�7�Zѳ��1�I���}��a6���j�����Հ��4[F�'*ȈTP�֓S3�����䟖j�-�Ut^���2����=�M̊=�fu-N_(L��ދY$X�����H'o.K3�Z_����A��h~��j�x �>"���x�����v�cnܬ����|�o�M5?�lU����-����E��l�2�?�3�y.��x�셯y�t�G�N��^�R|;�6�elx��8�j ~�z=r#�۝�����͑5E���>'l]���T�le�>&�VkM]�x_�1���c<�cǿ���o��D
h���rR��
t1 ў��S�}b�QCQ����KY�o�Ąj������[��&����6b�q|��g����k�Z_�.S��a�<	��8H�WW���|�T�o���o�� ��o0�'C��g\{S��7���$����]��`A��
����O���}IVB�=��T�p��wg���c��m�W��c��*��;{h���Pܒ��9-Q��+m�_	�����@N�����b\G:,��Y��4T��ˤAR��7�����l�S4���a���f���T�פy�m'o��_�*Q�Hi0�2j�ʘ �:�C3$�u��F�s)���c�h����Ȗ�E���S��mHJJ���;�����=!��O���&H������(aI��2���]ҩ,80�TGn-':��9���y�td�}�m���HT��5�1�R��J�������h��=	D_=s��K��5R�I��d��J�� ��) t���$����P:U��<P�#��ȂI�r��UU>(Dy��Q���h���@h����惦�o�oZ�s���G��(=���\WK�h"Pf
4���)�$��B�0	H�]9���*�%�� ����2Ȣ�K��:�h� ����+-T&����ӲB��~_��*������6���~L�7��PkIqE���]n�t��.%���)F�k���+k��uַGf=ͭ���8/OX<�*���SJ2!pF��_�`�"��з�����k�2��S���q�E�I��0���ɹ,��BU#�!��Ϟ���6�	����aP�E����ɑq0�!����RqC��J�|����8>Pqr�<�c����{�S�D<+[��ÞSq�^g�_k�"�|}E�{dђ�0a3��H�z9%�(�\��Bn >*��5v���?h> 4UY�����?�|���*���!�GpU�����9[t�vw��m�6Ac���g5'���_�2��F؄�
���h���oP��e�����_,-QU-ۊG�a�]־^vb���,��h�?B�SJ�'B5`�L�.�W���FW�ğd�|uٳ�� �z�
>z����c��<�9a�>m�77��4kT1RXpw]nMR����mR���:����О�
�g@�٪*�W.�Q�%�WQ��mf�ݹ)Z�͖�G�3�(����u�
�I
e7D�;�뢕�(���)@鬱����#��c�GCg"�rg��(E&tȓh���^��1��ʏͱ��N� E�=&*ʧ'pi��Qa 2�zm�UIҍ�x��ZL_+�Oc��ՕWG�U@�a�n�{��-�C����(r��^�0�D��$U��$%�RIe�����������v���g*�ƹ[Q<�{��0�ܚ�����s=������ ٸ��N����M��ի,�sT+,,u�Au������0��멂�I���tHӺ8�y�{ݯ��Uz�İ�A���7�;��g<ۉ���O���LWȬ�q�,���)��ggEN~]_s֦6Z��7,͛mY���b��U[�*)!�)������*[D6�ݢ&Z�'�ݙ�v`k>l��x`	-��|d��H�}DC4¿�9v����X�B�(�BbǷ���$D;�<_��8O��C	%�����l7���N�v�������v����˧Җ�e��9�V�aB
}!�)�]�𕕮�#����٬�Q�.�ϡW�fp��/y�N햸�j�����9e��C���#Ʊ��R�#o�l\v��#[���[��J0��?�;$}��"nd�e���=FAi�>z{�M�Ÿ�\jrb�m��h�
[VyUg��+�{�������H�`I� ��ո5&�E����߆+I@a��~�7Y*�Z �]Ĭ���3מW� ���������g�� 0g��u=��~'��r�^"�
�s���;WuCZ���V��a�� ����b1an�+�y�1�^�D��#8�|Y����_�t��ww����aѠ��;	��	�N���	��������^}��޿������g�鞞�1k�k�3��J�I��D�'����X�Uk.��*�@i���{����$Od��^�Lu��4�O'��o��Ȁ�x���Q1���|�QC�}"�Վ�v����{A+Y�N�S���!Չ�Y3��?���!K{L��qo
�DN~��4+��C�=F �,s�lњI:l5!ǟ���KCX�i�{���,̋*���M���A�����[�2%\\��5+��O�T��Z�xr���!����l?�<b�`#���&X������J�-
���^� O��S�F�Ll%��`�e(��e{���E
l�@�0ͱ̋�ס)gUEH>/!�ҌPVޫ�p��u�H.:�z=��i5�%�ڜ�.VQ�B�|S�A�(�����S��ŝ�ߔ�]{���n�\C#��iu����D�ƕ3n`%�V�*b��̗�yIx惻��Q�>�����S��������b:
�iɢ=.<KG*eEEs�S�^��J��#�A��Q��_*��DS�M8������/�7����_��$e�4����$���������o����C��?ߟ.3g��:��w�,�YU#2�d|�z6��\G��gLtW��dև�l���zn��-�P?�݀���S���S�&��҄s�D���$H0cC�܃�+�_w�X��>?��Eul���њ�
}��E�S�WVԶ�� zKW��[�@�%3޿]�&�ϰ�wP;�_˶D���X��M�#x8�r����m��ZŌ�#��Q�"3�b�r�ާzF{O�c~"ę���>��ՙ>�n�	<8���{:��h瑙�8~^J;�l�sךZx�WE��D�ma�$5X�ui�qhD��$FEu�+�4Uڜ1������P���N3�Dr�t���ڋ�ZMj��̤&Y�з�������1D�LR�:R��Z8F2�Q��N$KT�%���_���,��@��B�7����9KQ�kmb՟aE���\b�C{���JTF��U���A-J��0zQdCg�/�9s(�#f%�D�w%&�C�^�x���ʊю�y�4n}SэW���7vBa]'ըYK=Ɨ���0ͼ�����+� A|���B*H�4U�J�n<��QZ���n]�-M ߷s�iF�8ÌGƜ+x�g���n!�'����rzĞ�b)�8a��� ����ͽj���9��h����%�mH���lҘ���7ce���"Nr���	;�F�gE���C]�A�`0O��4���c��J&3��o�+��Ko�*��2]
�	�v��Z��&7�p�-G"5���˖8���5T��l����&���#��e`e�������Dr��9�!��3Y��*^��,R8�D
`6 �CgD���*�#gj��2���]ϋ�:�x�X?�#�ɰ
�8?������OB��$k�L;���!I�����S��a� 7��j��� ֊�
ʩ �~����;A(��SA���>^���|��JrGn�w=c)n'�x��d��`�~����&����+���N�$����J$
2?�ଗ��B�s(�F���+|\�wD'u�$]%^���,���ŢF��N��я������b��Xh	�O���j.@h�-��/�ۼ8�!�~��b�P�	Bu-�D���� �/仹 {��T/h��]�K�	+1J��\�=��N^���	L��O��)�~%M�vΛ�4v��p�#�Q-�N��ٴ���2P
���O!SL ��w{�dP�r����s���tJ��7��GqO�.�0�f�s~`�s���f�����Q2�Wd-���m����Ї ⲹ'��� � `���5����y[���9��ΛO0QgΥߴn�$�,9�A~�9��-�Ķ+u��/^v��~N*I1q���)}����ͥ�v�6�p������0GL�_v>h�j��F��:{��>h$1%�����<t�e���<�e�~�����ɴ�?��X|��Q�Tv�����dG�Av�b	Zʝ�Gr�d`0�����a'ѝ碃�{}H�l���E�X�γ�Ӟ��v�tl����fV[Xϔ����7�F�rp G��c�Y�	���֞���@�fud�)�ߩyC���{����0�Ѥ�����ޞC����"e~��_�O���l�׆񰕄*��B�Bz8�	�V��ی [i�X��n�/L1�QsW�:9[��yy���
��/�_��~�v�$X]g��ӏ�w> �e�o�|@YN��ӝf���@S���HF����fp��[�C+���J����
��`�]�w]�1�����BW�G�J��-��ݚ���"�J��̦�$p>L��M���6�����!����Xe
Ͳ����u��=>��|�+�U�o������.��H��_;���s6x�9M3�@g��$�}/J��LD%�:.��h&=��f��)k�:&]X��]!�j�U�1�=�+崂9{�ɚ>����6C��N5����l�� �M��)u�Fj�W���:,/�B�J�����k����o��ɛ0ͷ:���$�`0�=����Im}#����ΐ��"�aҍhJ��o�M�^X��h�l�����=m'E]R�Hbs���#�����6���[��4��χ�*�83�Ӆ�-%-ć���<�WOf�P�խ����RŶfJ���E��e2m�$�c<���
��m.���!����0��Y��e6����>j���zl�q~(�)��)J)W�����%�:� ��iW����s��K�,��T-H�?��+���"����LW5 �_��	�˰���͊`}>�Y�Qf�#��I^����B��JcE�c�gV,�K�^�~����r�fv�'9��T���δ���A)>��d	#r#�[��of�D�����K�v�L�6l�M�(k��Hx>�ŏ�ʏ��;d��ʫ�a����Ys�X���qP�>S#��>,�T7�~�檫iÒ�ii���B^�8T���]�2Ԙ��Tú�R^�ݳp�$�+ю=&^����VMe�q��ӯ�~��Dlp!� �#g���Ԓ͟`8�y�5nq���K��%j=���Ѕ���rN�c�z�����5��b�y���ِG�M�ՙj�����Ű��@�#rE�%'?�@ue��2�7���*��/8v3xw�plM{�-��&P���&rǑ��潹���)����H��:����z�E@|$���M�Q��&��J�X�\+��+�����7)�<b�׋q����/�}"�dTq4��H�F�l) �N������)��K������|�L�FAL����!��4�2[��g+<��ΙO˙�u�}��ݍ=�/�WG��w� ���ʚ�zf�vvu(����*�O�p��M���t5 �;
�@�����wQ_'l��mǁ߻ �_�_~��Ǜ��ZkX	g�h�߯�ai5��Vxq�G]^[�e�%HcfÄ�/�:��|�p3lDǬ8� 0IqW�Ǯ�I�K}7$��C9���������p"z� ��᪉� �n�D����������#/�&aZ��[�S�D�Nem���1���='�	���v�x)0\*��8O@�	<8��rRV�~��$�<Z�b��,����[�wg��$�	�+�b��{ �����0Z��5^�JH���f�=+ۭ�#"
<!n�D�?�kч��rB;��A[7�7����B��N;N�T���ݐ#������e5�P������1H��fI����N�����|�m����	A`X�R"SZ��j���a�I���?�<��	1������䲂'��d�'I3��K��r�=�:p2Oq!镃��<h��b��E\ƹA��Nv|0@�:4ϳMK��
�Ae֦�|����u)�i�����Q���}M>�k���n?d}s��e��]7�(�|����ոk��Q 
�jE�!j��D�B�����F��
ׅ���������(�c�>Y��>�h_w�9)�eUN� >�D��8��VJE��] "����zs�\^5x�����
Α�w�p+Ɨ;ĺ����Ӝ�����`���xYadɞ���� V���Pχp!��q��6 �Y������c�p��q|U��8@a�N�-�"��ET�a`~\��9�G4wK�JQ���4�|���Q�K<���{;K�s~�{���cI+��)�s���M�^��d��YK�����G��.`V��`�y�>��)�,�.9�۬u�1�nsT\����������ֵ���M'�t��,�H�#��G�o�m��x6�?jB��*����t��&�ID��Ib�P�y�Ot �X�b��3�#ܲ�|�Jx ɸ�lΈ��su��X�,���������5��h�F���&)K��J`t�f��s�j2�r�Z�{Nt��@7V��U�e��G��j�(_�\q�n݆|.L�ܱ�U�&��U��B��)�]��(T����R�w'=r���,D4f�w~��q��X��|+��;���E����ۣxp��)��������z�D�U
�3�еCQ�}�5zɞ���L��y�����늓���>䐮F�/P��P<���{��0x�Ʃ�$��bW��65�N�������8��!�ޓ����7an� ��q3t�$ex��m���Cͥ�K��~��~(��
%=���	�auH V5I�r�VY �#6׮<w$0}�hq&a��Ir���A�B��� ]:(j.Z�"��MV��\�-�ԉ��+�����k�=��K/�N\Âj'��i�K��a���j�����y2%�4��'`���\>�޶`>��cWNGMnѕ
�ܕw���Y��'�m�Y�Y�@Ҵ3JM��_<�I��T{����N��n;IT�ɦ�HQ�D+;�u�jM\ŐE�[+���T�YEq23�1�(]2|Ξ�w���@n<�3=�\G�nb3�ۖ�o���lig��*��,�ل��|��ڶ��=��,j�S�o��w
K�y"U��t�+�긏���n58K�5�cx��[阫`;rs�;����͘����e���i~���z�x�͌�2�M7�BVA���;Dp�'��~W�����X�[C(�׋�_/70�F��0��C�<�y9-���%�.��Ozj�q��d؜��O�Ӫ�����P�V4���#0�-�����Q߬��z��@c��	�$�K0����NY%9`u�R����]YK����s�;������J.�/P�N��V5��PI	��Y��/4���Xh��y��-�)pv��M�nκ��=���. �g������W��;� ���X�YZ��1�T��V�q���#"bgiB�3���9i�xMg����,=����f��y�� L9ع𩜲�\x�r��wl���e#�FWlw�w�-�5��^�+��U76H�
U���HQ�E���HvBM�$W+�2�۞.k���X�R�j($�P �Bm,�YL(!ެ�.�ҷ�'D}�:�yE�W�#q 
�8��jԆb��W�	.J�ދ���"�@���%:V�L5'b����&M��d�ߵ����
j	1-A	�����/Y>�W�L���؋��!:�y<�p��8�.�Ŀ�>�3��$A�]�t���~5�-2c ���VhCO�20��G��[S�F�kz$�yz��:xm�8�JHJ�����Q401譍���0�O���w���?/��A�蟀��V��/!���B5x�.�ې��F��]o@�!)2ĵ���^F�"#����ǒ��orM��'!OQK�J���=�x�w1��������?��A����[�E�ЦX��1G������?���`�d;e��Z3���Ͽ��/��8w	%0�o��l���2a�'wW����,�R������ݝ��˳�$

ʊ���F;a��(~'�3��W�
������im�_o�5SY4�����f�|^l�ITH��p��=���@3ok��c�Zz��6���X��-���˽P����1�D�a���� ���%���Εa�|���pk֯�tk�)m^(? �iF��&��*�cP%x���$U��Mg��%Pl�C�2{!%�b�|�2�OARr�::��(�ͣ�ﶙa����{�t���+����D�?j��� m�8o�����q:�̌��PC1��HS��w?4�~�+����� O�v0J��3v����]�໫��s�����Dkܘ��Ǵ۝\#e[k����ۇD�m��mA]�%J�x�5�iW���ۧ�X��������㺯0�J\�鎙b;�HH���<�����e�|�ܑO�1������b���^lw��L��?}*�g}|i�xݑa�{����eI�Tv.�MT�:'��3H����������._�+xd������y�޵�&PÍ�L�n���e`M����Fhr!���R���0L�D@�����z%��a򞊐���h����Ƥ�:NT��G[�U]��b�E���@y֥�C�,�K�.��>�����y�ӥ$��'6̠��<����Lu�ZH!�h���?8G�Ew�h!�
~#�����**�;��2N���--��
_p�x� �m�"���fc:���DTo��JMf�z�]k]�a�L�X�I�P'�	F4�r��ɀ)�ROڝ.GdW�,Zl�Y��
f�Ac�ړ$�>��u�<�Qh���\��]K>���1��oϢ2]��8����-X|D����'NW}~�R;y0T�{��a��*�JGZ�QB��d]�h"@�2U���cJ�d	���r�
 �p�S�T�?�1����.�9F��NѼ����=�8��uLy��3�{j
��Ҿ�IL���d���|m8z�+������>b2�&L�; +�?p��60�J����D�@�t���ګ}2���aJ�b��e!� $�u�F� wmn�~;�&I��oL�}�;$,N�Ծ�uX�6H�"ϙ��˥E��n�Z�>!f-[�"5
V!,�"1��GS��ό����b� 9X��+��ީJ���yY�y�5�����̋�Z����D��q�|����O��'L�J
���N��� e�!����5fʓp����T oXN�;�̸;��PZĲr��
x6�����Ĉ�v_s+�
���#�P��߃q&9!�j[�� a4��I%|��C�@Q�=�[�4���bC��!U��x�T���Ǯ�U��:^�?n}���ߗ[�2<������V����RĦG���K�n�rU��⅙�.D�ENf�[C��*�}��Iƴ/��D�N��9�]��t��~z8�H�Bw����~.�q�"(������܋�O`�&�8�L�>�H�``�z(������������N���W�f��u��nc�4��g�1�}*�A�@e�]����VWN)�M��`�p�r�{�V��B�U�*܁-����C��V<��!�Yn�A�� ����!Yb�=�"	EDW�}u�� f��N�a�w��(ta;9�8�b<y�EE3�+�c�@^�Q<=��P��'�+;pA~�E^�B��{s<P�����s��p�����1�Ѷ�8j��z�$��zX��y�=��K��ox�տ��(,�5y���z�f��(���G9O�Q�۹=�|6O��;|���f�zvg9;��I����]������ �����Ҩ�S�M{��U\1�|��:��&K���Kq�^���i�P!b`'�E�[��������l��k�♌RxY�x�o5bFk3��Ӯ��d=�fQw�u���g�k�4���\63E���u��Nȅyn�A�av���4s�Cup�}�o�r��7��Q���d��_!Jͪ��\&��<l<ۅ����V-|��Z@��;+�`���9a_I���k�Q�W��p��;Y5���[�68����_{��!���@\���}����oY����v}�û����8T�-��<r=݋��7n��[���/�Z���㎱	�CU1���-��2�^�m��/h�m6앲��-��z�k.����t����⠏[q�%���پ�e��	0�i�����ul@b���V��l&�����8Dt.����UQAgŤnR{s����\�>���[ߔmD�l�j�Ov_�{�j��z��d�۳�Y������9{~�H�:������?����A�?^Y����t`QQz>���J�)fI}��kq�	�9�f,��\ޱ�e���Y�9J:�����{@On�kz�H���:q�q�L�������&k��}���6HP���h��b�0ث��ʄ��;U݀��6zvH�}4����qpf�[���A|NĴ����V��|ڂ)��n�6�/��K��>9�45"��� ��	��b:��M�!�>Op�0��4l��B�ֿ4���~�ݺ��)�>)u���t�˺��4Y�����evZ�-�x��g���ݹ��#!O��?����'gSU�0�FQ��=c}�j��)3s����R��zj/�}#"�#=A����2(Q�.���������&�Z]�^ߒߴ�-���0��껨� '��qz��VO�l3Ի�e~b��a�{�hH��(��"!�؟@�z���M��^��y��y��7'5w����V�"Z���X���M���xn����z�VvUm��{�W"���r�L�%�&�����7�9Y�}��5����T(��%��n���)R�TTl�F�{d�lk�2@����QD}'�ZU�ϸ=�	���8�e�pF�j���k��^#�*'܋7�6�m0)�9�P���H�p�D��H��h��y�ePc_�O|��z��1)�F-Z�j��)ӡ-��Fe�Tw��Ѓ턛�$C��G�K�_�����{����E����ǲ��1q��M41��*耆�>��? ��,�z�"��ޝ�T�~un�{Y�
�KϜg &N�*���mת|'p�h;���рɥu��˒�6uR��Jjn�/^�D��W�6��N��~&7��#XE���<�r����O�����^��]d��Oy6J{&n��}^'&�~�N�Ef�2n��!o�M�~"|I�dyP�䚒;6��# ����
7M�
;|t)=��C&!�R߄���Tli��bk!|��j�o�$��C�eG��O�C}���x�͎8Ň���m�{86~�)n��l�_��<��0�N�F�����}/K��AD���Wl�C���Av�1-�N!ͯ0��t���J5M�I�pD�U:N����Q!Q����8��/���s�?\G��\��7v�SS#I�,Z�6v���T�%��y�]xeV�vf��?��Vݣ.��5r��.�I�}2!P��V�A|Z��hj����>$����0��6.;d��>�4�e�����LZﯜ2~�G�Zش	R�ҳD"zHHxG��I���a@�7g9� ���30�+�s}𯂻�r��3[}�g[�Q�@:�J�K��� ����"�"����D (*�F#�hl��x�&I�tY�^�]�h�����8y{����˯gR��sd��k(�����il)��ہ�g�ӶŠFo���n#��Յ�0Z�<����c�9�=�`���N;�� Ҁ�XK���KA[�7�^l�s�s���hM��a��5b��+��#EUҪ�k��Ib�j��d�ɞ9?����x��%�$�&y��uzh1��Y����>�,Ϫ�É쎘	Ʈ���J�M��?�����|�����XQ���'��f�΢���*�^�`�P�	��M�a>ռ%�C9N���4�e������Q5�$�s�uc�=�Y���2�$�L��Q���1���9�m��ױv���Z���[?$a�\
_MLM1߾RNV�zW��L?�zG����w�<�-�:���TjC��,J���Os���`�8��6*~�t��}s�����W���b����R�\gUb����ij�����+k�]vD�t� V>M�>�]�Gв�Gg�Q���$Fa�Um+�l��)�m��t���������	�:�Ek��5P',: ���6��[���Xߑ��1�7Z�
���蛂y}�@��[�#Q��c���a�׊���V����F(&d������Z�`�?��}�5��x�ڴ�߫GC�fO��d`'��c�D�����wj���H�T�t42��sHk���U�U[�e>_\��V�)rt2���U��sE��.,_�w��������ֈ'M�H�>�SS�������9Xv<Ϣ(��i��V�p�a�Tc��C��m���X�}�C>�Yun�IÐ�v����hR-Q���P���e>ʗ5�x~��>3��<�!�Jk��Z��݆�����x��a۲-~�}v�)�Q�{���F�+:��0��a�[7����H�{��W2��~<ew��h�J�O���C#�s��ֳ�X�r�WVC�^�d��MS�ZQ�:$�+.�(�d��qp+v7����D�/m��5������{8��_�gZ+��̋rk��n 0�㉁K�^��徫�����^jz�Lj��"٘.T����Q#�+q�v��Jց	��?�Y&�|D��$��P�����W�s���J�8��z���WN��x�W��h�x̵+Ga%��Ҫћ�k��2V�$V$~������1�Y� a�A���k��I7���(FԍE-�VX�P�P#�&`Xl�MYx!t2Y��f9m�0H��%	�f{˶M�U.�7KN�KU�<�A���P�q)�(�h�gm��>V�񙜨�CŻ֚����6YS��dޭ+AO���K�G:�yPQQ?�,͌���z�#1�M!L��K)֐7T�}�1NKS���b/2.��7��Q��ػj8*r/�U����miV��@R'f��.#���+Ԁi����'&t�q��[!1���C�7������t�BV����B(AV	�&������2��^ࡗ4��Θ"�Z�ao����4}%��!z	K:��lNq��)�W'�>Ym_^�A�{�1v{+�0[pl7���������H3�\�0}�ƍ�cMs;�>����.�x7=8��O,��i�h~D��S���5�0��D�S�,T�0���~�㙽p�g��q�R`���0���Yv;ȻR����-r⃿�!�K*�f��!t�%�%k�a{�G��0ᄿ�m�S�!H1��Z�L2���7�;AJ5{#Dx�3�Y�F�v�MZ�f�&N���l��C2n�{����eѨ�PGG��s�E��'�;J�}�T���a��A�
u�Y)HU
t�'d�!$��S��6}�А�r�������T�k�͐Ő�l����T�ښ���ѷ�[��a��ڧB��;�؊ݶ ����N*��;���~��85�*��1S:��Gr�Vf��sC&����G$��qcvl��a���|m$�zS�x!//5���jh�����a$�08���ƼLn�
#��Gg��lc�4�Gz��u=v�7 S�*�����=�0�Q����P��)�����5~��w�caZ�x��ņF�ߩI(B��2��I"�٭1���:E��N �sc�h�9�|ۂ6sX�VDY�Sk�N�� 2X�@E@x��Nt�A�Ͽ�M�R�}M���_.�PK�f�Jx�Rϵ����%��LPw�(��
l��-���QY~.��1����\�GYN^RӀz�R4��(�K������|N�L�-�>��gy<v�+>��������~6���z΋��ǩ���ysXpjFOp��Nq���F�*�:1�3��i�ʆѧ�����)aC����Z_�����K�!��u���~�xE{��/Z�+t��d?�OGP[l��N���/Pi���貁O��Ǆs���Dj�}-|h�g.*�~� �.Ww�3��ط������[S.qJ�X�g�9�6ʸ�}{C�w�c�737:�Γ��5ikL� 17.8��u< ������	����w��T���*F"�='�~ZN�{z�e	a<����g:�<W$�~�'�f�u��5-�YsxW||<��	EX��c�F�-B�QU���B0�ϊď��H�����[���ݐ�ŨFQ�]_���F���g��� b����F~�DP_>�FGa�2ȡb0$��@��( ᣯ9�όoJ�������Jͼ�4t\�V[����J�(tw'zЏ|Q��,��5���� ���Ɩ��-�r������E]�.'�}�3��cQ؃��`��P�R�	��%��*r�mQn�gn�'i���مW���y�;E�Ͻ����F�곦�Gҋ�q�m&gD����T>d�[IHZQJ��L>�QR��4���LN~�������%z��& ��G�ǈܷ�����~�	۰:�%TGѰў��I�0��%�Wgx�ne:S�σ��D�ڮƕ�l@Zj�A������7ǀ��~�s�2�w*C�ZG��>!��r��Ɲ��h I20	e����Ks��,o9!EVs�&��0�F��,�U�/S����@ٷ�Y������&49�w����<]� ��:���Vcg��כ�L�t)�ؚ��+C�%��mo G�)�Ax3�-*�:�9$P��ęP�P�V�"p��	�+g�OکF�~�F�%����~=>�[Y�%%h4�-χ��߿׻x�>7�dd�K���/�`\�9Ț����"`�_PE��i�6��ҷ$�@���/�>r;JX���5�Җ�Y�֘{�*�Y�♫��� ^[��Z���=��f��~��//�[ɛ�}�+���df��t�U
B��bi���:w��ȇ��|#ղ��ww����L�جYC�>z�`q/������^�������n�g��U�	�� D�֐��,X����{~���N,��{B�~�ٹm���˜+����dxsur�&��\U�V!�Y��
y��Ր��4���)i�7,jќu��x�|^p�[�#:-t��P��6峷��P��k�\5������>�O�x� ��#�������}��	�_ ��� :_��k�¬�ە�h�w=U�(�Nc;/+�m����y�WDp��>�)���j���p{Ax ��������H8ֳ�g�}����3�S�!��*�&@?�J���er����Ӥ�[Ox��!��;X�7R��*a�u�>J��>�F)�����f޾Z'�"��~	��>�pn���f��6����I���9�=ۙ�HF�"�c��R.U����@��>�a��P���N���9�V3��~�1��J��N�^��H`R���ux���(q��g�^���8��+q�S�+r�,�v�A>50�?�l�u~��qZ�̞ŗ��g���vR�
fZl�k�[�Qi���Qf��g��&���և�hc�W�I���0�1/d"�N�c�T$g�D��W��a��%l�����J���a��	m*/�f�QnRu�1�lU�61���-�cYs!Y�Y�N9[&j�ͥ,Z��#�7������H! �&�h~g��Z�/��M�'`>���2Du��D�
�WT!"���<��+���u��]��lQA3�
E��g	gŸ���3�����HPg�j� ���<}�$�7�h'��_>��ۋ� �\����%E�ְedSY��0g{T��;�Ҷ����dE��2o_��dk���x;�!�*=~�hj0�!��t2b�n��"�����교ݔ@I�R���@�!�J�[挶�.8P�eS �B���]LŌ���#5�r�+"j�v����ؾ�Gҡ-`fp��b��6U/�jOǲі���6P�_�O��ӻP�K���S���Ȼ�#@t9Բ8B����!����e�Lݺ=x��	i`�q+��p�Lq �\�G$��<q�Q�ؿN��ҪXV�3�4mAm���\��V�zUk~�ֿv����ڣ�#�^�#��F�,j1b�U��
���j�s���F��ㅛ��$]=�c\el�V�u�J��$�v]�7�?Z������ _�=Z��T9����Ih::���3� ��G�77�:)e�;l������6Y6vD��_�Ë��]�,�d5(�DW�����J/o��o�ܝ":Ʒ��'��&��v�+Zf��<謣��I��5h.�_�^6-L�\_�&���<-+p�$�j<�Is��p�2i����?�{^�eT�J�~��N[��{��wA�;)"�3��]
���b���>�����w����h�H�Z��6	*�^�1�Ç�������`�	�Q~���2�@,��lB�|���@�F����������w��J�-mCn�}����7��)-$ẉ0�*���6y�.��E­;p�M�·۹W5�4�0�I���B���f^��,Ÿ(� )8�ԾS/#:���w�J|u%;�M�	TcQY#L�7��O���թ�̡���)�&u�I��.5#��"�bT��^.J#��N��y$,xݼ/�7L��+�W[U�jp4����2�j7INΉ�E�������o����惑9?<�I��R�k[��o���P��ݺM���*ĳT���h��7��,�̤'O�n`Dd��@_O7�N�ld�{6:����O�|���]B��5���i�eB��@�K|��%;x�5�(c2[� ��sj4"���7;O_?��R�!��ƭ�dh5�/���q�~��*$3Lu_�u��0���7~&������ �犸������z��&�x�^�
l�C_N%7��1�<�=Қ��~����w"�:�����m���&��N'���^�xF㴐��j;�z}���7(ӓ�MeP?T�1�;�W��OU?��Q�0��V/�F�K��=�������Xx܏r-�a� х��3������$X��e��!b�6�_w�j�{�*'���'&1�c����I	}^��ڝ=�H16=�>e<+O���d"#5�ޮ&L��A�B�CῨ�ݚq���":�\j��e����ǘ�yV�sj��p�$���)����_��P���h�υ_�G7�A?�]���tYPC�B۬�
�qH��җ�Z|o��Ąm��������¹��o ���A�oe�5�N���oI$�Bm���l���E�A�J����-�f��Ԯbz�ae���1$af=�&7Z/�,`��B#@���m�nG-'6K�s|��ց�>��ҼN�*9k�I�c(GF�f�26L�$��|��(�4�f�9h������TxPB��հ)��ҭ�^�a}\��⹛dSyy����r�f�g�p��Y�9���(�K�6�8P�FR؎�x_�a\�X��}�yQt*������
G��o�F2D��o*ɾ.�Lw�)~6��)��:h<#�U�
�u��Փ����5<�󉨳aQ��.�_~�,m���-�=�2��Μ��� x�I%�*�O�XhQ�q�5���&~�(�����0$\M:m�m�:!X�������+�X�%�4v�A�ǣ��Y���l��7����o�qmr�2c_�-�:~�qO�dj_����O�`ܼ�&A��T��%�K�&���� � �`E/�#VB����e�KH4�tg��\w���	K�P+#���z_�l�Up0�����ڧ�z�Z%x�I�n�]�⼾�1h��Ek�����*~.�K6�y~�K��e��i͊���R$U���۳lY��U?<:Wk��#YwoаMz�<��Ņ-�OL�Hf3�V���X�y�7@��
ŭ|��nz�A��=u�T�_�$�� ��d�{��Z�]�M�%y���jm��z 2qh�|���J@=EC�n�{�޶34 6'u�S�$By�6L�l	T���U��� }�6yx�l���&�><��BI���2�}��J^b^�
��M��b�e��Ebk�o��2��]�қ�aSd	#�ʙ�l�X>Q!2[�>�#�$�>���ӊt�l�/�I���>���k��p���}"�4,�Z�\�O
��ּ��&fWeD�]��_�!�ǭE�ó���}�G�渫:Vx�!��9=���o2gYRݻ�5�_d��牑�������EݙS��ru�	�΋^����eQ% n3x�nz+�M��U�P�eL��yQ5:'�x%װ��ϟ	?�s�T�?V�3�k\x��޵?��)�Dh��/!�_q)恇��vvC��?�*J^@Z&�;�ܵ&[���v)��������)��2)b���7(���!,H&�t8^�q4|xɱ��=A2����/��Đp#��M-�W�m��P��`{cVZ8P�N�� �0e�zѪ�KԳS&���p*�6�9ui��m`X��y�{�h\���#�f����檨p%��vH���@r�,+�-���Ygւ���dM"�y�P`��)��(6G*�P�!��u���/Ы(Ds�z����S[�����i�F ���	 Lb�J	5- Mx��@�2h��6�Y%���V�8�ǲ�`i\����v>�_�/kd��<�(0g��I�א���������ͼSh�/�z�8z.ω�Q歄f�3Pe�V��[�wc����1�J���L�Cs�[c��������"�[:h���dT��H�38��@�vKl�9A�9���@�{?dZZ���,���iT�.8텴{C�X�_^S����Ĺ�F\��4��(��?B}QB1��e��XR�#t�+�v�v��v�G��Z�ɟ�8Z�;)��,@�p���Nzu� ���{Bڒ)q
��%O��b�d��_{o��	�w�tY����>�/>s� ��'��}*��pH���hY�c����r�7�x\5z�g�aM��/�����(��Ľ��hƿ��Wx���'�H��������N,o��hs���j�_�(�Yt�0E�z�D�I��i%�)<��5D�5
�VN��Ȑ&Op�ڔ�!Mvh��h�����^����^��cI�8-]a\�W�����Q|~ɂ�!i5�C"h�Y�#@T_C����B<^`8�s��B�i����� ���݀�xTN�&9m4A��"�_݋D��O:Է���,�2��D��z8�i�H�`A[`��-7��9�~m� m]�֐�h:h��go��`@����崋�������W�&c��\�m�V��pL��"�m�� m�����jK�x|=ySH_4�A[(��(3��I����Z�\H��ᨁ�s�Y��s�(6]����I�GW.@[��!�� L�a���7���A�ǳ�i�L���E��n��K
���!<5�Ƭ�@��v����\��+���6�L�#�ql�8��0���o��]��)/���Ym�� -:��q�����1�6��}4XЮ)���*,+r[;��Nj� ��t�7��k�7�ӊ{�5ZMV��/��o����#R���_~ ��W>��ΕO��J
MW}α+�R�����~�\��GqU�-#�6��Q��;4��TNܴ�\kh�14
�Y�ƺ25,6'��C'.���qw�N�`����ل�wm��ւo�D'���pN��`�ϕ툫�����Q\��*�i�Gˀ#Z�Lb����G�n�C	5%
�E�(��`$#k���m%����A�@Nz<r�h{����	(���i!�����_#8mS�J	#ν.��N�n���8#��)_����d��������6��J4�~�2���MP&ȞO�i�=)8m����Z�ж$,�6��5���Y�S��Qa=�l��x�
��<�]'�+ٛ]�<�ԭ���N�N���L;'��-i(L�Ld�g@�{�����A�.�)�:(�I�j~z������_=z\�6�����-	˄xL���5��פ���aTd)8�U31�R2N��|�
_�LG�%%���w�F$h+˜h7Z�x���8a�XtT��~�8�B�!gYZ|~�brZ�����v{�
?fb�\��8:���9���z���t�[>���@1�ʡ����ywY�F��{bR㙴'�ލ�*|���ꊹ3q3�����={�o�5���M9�X�L��R���w��ԧuN`��kL�J��D�l'��y3�9e�94#��%�u�C��*G�LE7t�1f˞������n��5}d�59����i��{!6o\'����_�ǹ��o|�� a)��Wb7��/�	�_1�=_�t��<@��|�4��E��P��r)�W:^��#˵S*<L�b�_�̙ҕҿ��3j��oܸ����E�}ƌK}q3�Y��ĶJ��'�"E����8���6� �1��\B���
�)��gs��F'ڇ0��x�	C�#���K/�b��:�X��ǼL���v|X7P�Y��e�&���k1
ܮ�3���ub���\
��܉���(p�R j�����;_�K���j=�]`�}7뱖f��^h����9����)�����\��Ɠ���G�����5¨Ȓ�R��5z����8�\\�Y�}��X�Ů�ZǬ������oO��l�n�޷}-�k� -���żQµ�1�6\��E��y�]�cV��O_�[��%����������*��
͓=�y�@�@�z<iwKNyf6��ǳ1ʋӝ�l���L����6����@�������8;)T��C�cL�������=��-�^?'f=�VY�7�@+�X��5�ig��s��1��Օ��WL���k�NO�:߲1F�X�����6f=����Z����+�Q��������,�%�� �D6ƃcx;V5O��hou�F$�Щ��ͨ3�X�d���4fFǜ�ɻ��1(���:<�L+�i��� >�����^20NM�����{ /?��p�x�9jU���
$������N�La��`g�~C�v�ڇ��i�t��(��Z��y������m8p]�na��Q��4`�f��̇�4>�9*��h�9P�6���#��H�*��]����q�B,�.S��ncX��j�T�^�)�����5��&�����/S��&�I��:�k���{c��0��L%�\�U����ϙ��Y��T
�q_�?ܩ&�;gF�@h�9fm��V�P��=}2�z�;g��z�g�ڵX#�K��W�ﱋ�� �q�@�!���:'%��P���k]ѿ
8�Z\3���H��Q]���)�X���Ý�rc�M��ݚ���l�Z�ȅ��:;�&�Q�؍4��uu&�n4����}hi���z����~{�xoߘ&���tڐ�7���iC��1���T��jR1����E�ޚ<zU���O ����ֈ��� J��7Ͽ�ZK2�!���Q�ē�)`�/����&�Z�{��:|�W��i�>�E������|�\x�\0��;d�9�&��wb$e��)��\ck�C>����*�v*��Բ^<;��]�Vɣ�˂�&V�/�N��
�����F����6�c���7��c=�V��m���F���҇CW��:��nBA;t��fm� �>y��w��ckl����en�ɸ�۸ōu�$|�M��NN�d�.�(~��7hSW�����!�М�i��Ʌ��&�,R�=�_���$��*�Al�x�m�1]� �\�8}��j���4���vo�t�U���')H�ˬ������8s��1S׈���I!�wNZ�	Z�p�cFjl�M/-}������E�I/�����n���S�����&g�[�o��U�*�軖�H�bA/�.;l4H�_��Y<�S�H['�kW%���9�i�hi$"h�F��\�P�!�R֢e�c�c>@���gl�5��9��,��`�]�g$y���E�6��k��,}>�H� ��P�L!,g"Q3D��i#�#�i5�A�YRG.���1�X����r�HX%9����~�WI��d�{+vN4��5�WNY.�eդ���#��{���c��o��PΓ+~�T��|-�����Ռ�b��dm�́#��V����8�x���-�V\OZG��?o8-o�T*TJ�'�v��}�����bAK1�W3$�p�PN�8$�V�e�K����`0m��aoɾ����>�o(LV\�D��?ot��4v,�FaF<�����Cuc�*,)NƪiH�W�oĂS���9
��=Z�@�A���,���~��g	0i��W�J�.���cאa�6^Pjr\~3�R���h�'�ݒ���Qɶ.d�]��64�6}��+G_|,M��ZK3���\vw�'����N�F�q5��%%|��.��z�sy���j�M6���q�~@І�ٷ/���;K�Ⱥ�	ח��8_���&��E�z\����2;�S�"��f�O�M����m�^Q�eR��۰:��'�Z��N�g;�8ܤ�A${���V8��܎$��)�^�I�j�:��m3���[��Vf�������6�CMt��1/8-���ݷ ?���~ۂ�s&�kQ�s�g�VᅻJ��pֶ��4;��aߥ^���h���F�Ӯ*V�{�t`����D�O���%��	
1��K�|}�"bV�w����h��u:�n��I����<���ډ&�XV^������_>Q-���e�>?Y0��5y���\�������4,@�=Z�����������Y�@���@U�
�	�=��6'���e�Xd|nu�
%�����8f��A[���ҩ}�v����n;z������Z��k�XD.�5�r����:�0ȅp:�ғ4��I��_���A�͌5%��-S��^u��g"���w�)ǳw���w�4�hCY�س1
ȡ��/?�/���t]�K�g�ﭻ^���H-v��^������JIP�.)N�=v�u����������#�����(��;J������9Z9�"�wNS�:�=eF<{W5�lZ9��ٻ���_������P%��T����9��݁��2�[���.�ǯ�80�S�@��X����>��ކ��ɡ��?\�Wv��,�!�9U󼉰���Ǫ�Ηg�a0��h���+��������#.OE^"��(̌�_��]�4��c9�#�w.R`^X�ݢ��܎�^�>q`��������r����Ž+s���e�%���4�}��sq����f�
��qv��f`uy����-8R׏S�C00!���
�&ccu�����GL�����i#_���va�!Y�h9�p��2��U!N���l�q����	�G��cqq2>>ىK-�������/�T\������ppZ�_�V*��jǲla��s!���R�L�H4rǌ�'=�r�H�A�<�7Rs�B�y������m�F��0)��;f$�=�)��Gjr������TZ��c)��'\�����A���LZ��q(�IDz��R8��q�ǈ���A�M�kLo��r��%g\9}����O��r�K���1��]T���%)�6P�N�Ⱥ|��B��1�|��^���S���&#��W��qКm�Q�e�Ѻ~��7��:ڙ+�5�����F�����޻ 	��)B	�yI���m2X�V�BJ]4��z�O#�s�K�К<��kz��a�:�Ө���CU~Ƭv��h;�9҆���Sᘃ����O�<����}�yPKm��e�	i59m�@K�b=�~y��h�8��@�P`Cu���l���0=Q+��G-b����+f%k��]����"\��gg�p�yx
h��,��GQF~���h����X�s�
w��-�,���᫓�pr�����$�Z���,���c6|s�g�6�GIVJ��ρ�����${M��P����X	�Z�Q>[j2g��	T�%
_irD^9}r�S��c�ܹ$���j����O�q�~V/��t�p��Ӈ�g�����ᘃ\�..J�b!FLV������rx	�<~ro9���LLI�VR];�f��i�OrԪ�d��?���/�M&�3o����b�"a{N��x� ���]Y��7:��MNC��[zr�Z�̠��8K��Q]�L�S���]���=M�	/w�z����2���Lp���$���F��'�ʅ�Ͼ����"�Bݤ��1��-�>��B�'\��K��Ғd<�nY):<�>_x�}|�C8�ۦ�l\����ۄp���+��S5��u�Ξw�% 'E�͋2WZG�̤¦U)A	�j�^��|����5�7����$d����m@�Y��բZ�׌�us�%E)b1��C�\m�1��]�'�{�����~X�/κ�c��Fc]�um�)��[�/.><с�ܕ�[�q�Xn�h���(�I��p8ETXkߤ��[����e"",ܠ}hM>�c_N6�W��W����Jq�~p"ڌ<��8uP��7���w����ͽF\i��J��w��Wo���h�`�ZU��)h���F��(Q�� 8)9*�_�M�-}&\m'(����y��\ x����`���e�?���{ŧo�� 907̿�9%���k��g�T���]�����e�2>O�)%AZ:P�~��rt����NmR�����?P!���d���'����b�xW)�:؊��6�����#�u��u|{ɵ&l�U5���?v�>-Q#�_��h�N�}I���KJR�	�1`v=���E` E��y�@"g&���W�l��})�1v��U�����l�7	.J����2��?I@���\�y�����^�-��o/����y�1��z߯�7�߾��&�TB�{Y�7f7�g��<�:O���¢.���E4�ݻ*�iز(Kq�r���>����(/�i���������݇'�C]�?��V��o?��o�Oz��\���x|�H}����%3Y+@��u��b���V��ZN*�1}��3㱨0	+�R���<M���/�8ݠ�mӣ�c���̄R	㍈�IOm.�}�H��������P=7��9x��S��xu�~p"�sb���Ɏ)��!��Z�)�,}��l���ϙY/��Q*te)����JS#Z�y�o(���A�P�:U��|r�}z��l?�^
�Z!8"�}}_�o�N�?����V���o�<��p��>(օ�.�:�32��s��&Qm��cO"��ĩĈZN�5*T�'��Q��������Q�i�� �Co}i�xzK!~kS!h!n�3�r�K���Q�Ә�
��)���Ë������*���:��x��0�U���Ǫ��k���t�֟�����)�4+�l-B}�hX�c^�-*J���㑵y������J�;l���ljJAz���)���kN�!�A.�>�� ���J\l�n���4��h����'�Gi�XZ�"�⾽ԃ�����ɼ�i=7u)�T%�	�_�4�s�(Sl�)JFb�
���?�5B�8��EW~F�0<��$��x�J;� B�mzԐ�;�C-����	�X1���ӝ��T�88(��������,���A
P=�D�z̄���G	�?�5�@m��R� �q�cJL��|���*U8���w,�ĹC��ٺ�ta<�==m,�i���2줎���		M���/кM�$Fyn�б�km�Ɋ�G�@�2㱸�^���3}�{� n� ������w�И��w�AKN�K{6rC�h<6�&.����v� )�޽<�w�q���f�{��Ӊ-��w	��F�=��!�5�TCɏ���o+���eZ�_�mB�И8@�Pl'N\ľK=�����5��*H���V� 9���da��2�����擺��u]���K�ru~"�J�Щ�9�&F�\�R��5g��ȃJj�?2���QW��P� ���~�-M��u�n �oI�+Ј�f0O�=� ă{��T���Ls��0hg�؅�eF�F̑b���u�s�w:-9E���H%�R��2����$-���ϺET��ߦ��&���g(�ґ��ɂ)cY��r0�N�3-�Om.]�6��>ֆCW��2�ٸ�x7�d�	��e2h�u�⡮AQGe    IDATK�
�����P�XX��&����W�<��ab�I��=�Ń�n���5R�5�r��X�i_U��ؼ�YW��p4����� �n�FP�6*�;��O$8-�f�"��)J=���47�jq4��%
q��kt�A]����3]�P����*%�h��"]��5�!�\?�NZ��2���N\i���̢���7
�0x!\����+0Z�??�%�M�8ݒ�����/�O���7Y3�5�5����U���v�6�.�Qm��cޭ1-꺪ř���+��Yh ��u��>xR�/��n��ݬ���*E�m�3�HN�|^i�ԭ��Ǆ���<�C-��"��0E�W4�mY��;g3xB���N�?�(�����+gѩ�
��Q,���m��h�Y>Gpo�N���d��s��_�}w.,�����oo.��n���> ,����IK2��(���C�!�!�>^�ѡ���xII��?k[�'�h�,*Lk���i�Y�F�f�aB�w�7�[Zy���
U�5}�m��~r��\���e9
.Fs�	�&J -A��T�')�>��|�@�������*`�hE�qش0W���0fǑk�8p�Wlhnd9c���<����|ܷ2W ,�Bݽ�eDx���@����|d�h���í"ٞ�X$�����&��6w-ˁ�����p���3�Ⱥ<q����ӝ�w����)Wsr��~T��C��(�s�r��z���
E&D&h���exQ�{h����a�5}!yN�4�/s2N���*�㠭�K�����t�q,WBQ(]
�8/�A�}뚊t�q�^�܏���i^ʘ���kS��o^�!��奩�~�y��!i٥�-������W�{��9:Et��@})��Ol(�=�o�d�\���t	�#�A���-���xG���k⸻�f|�h�����i��T� -�s����íx�VtNV�sO��9XO����hn� \�`������8E=���=�SC>�D���\��;���X���%�\��Ƨ���� �2g��[��O.�M?<���}���C>_��-�|qyn"~gW��+���?_ݘx��ߗ��/�l�R�0otZ���_��Z�F��ǔzm8��i�S��Hlϫ$os��A��Aq>\\���u�i��n��.q)�z���V9���	J� R���a��߿o�E�sW�F���嵛/���y��Kݕ�m��Hq]�U
��d��?t�O�����G��I�<�(�ӥ��չ��KR���ο��~����緘-v�����F���P��tƦn��	Ը�)����0����8����/��s�ś��{cΣ�5<.���h��a���CW������ ���V��)B���7)}i�[�Z^C��9,\�f9:f�g����nq=7ݪ+g���t��q��,a�}}C�Ap�����)Ewf2�A��N�{ӭ�3�B�<|у����<W��z����n��s�8��J@@�>��8�??��mg�hC�3��t�Ը��2��ň��Va��g���CΜ���u뵡n^�p\w^{QLw�����x4���S]���`��JP����D��P ����\��T�ǖ�yx�����R$|�y 0��g��JU��/4҂M[E�7����m޴���xaG��%������"����S�g۶���w^������/�NKRx��4����nk+���=������b��G�A��ec���z�+ܠ�����|��$���BOPҷ�]���gYi� 5��1�\0��;�65�uG��<<PyG>��b��"t��]?A�F�i���@I���Tt �u�Px�Ql�cAL5����(���r�yc=�]=)C�X���?�.8�/���a����Z�����?o�lrǗ�ōA��>R[��cz����	� �{�G$(�F���8��:G;�O��9QM*w�E7�Z�,Do:��SY�61�h]U��!�Ɓ�:}�,���+�蘒-�ܞ�E�C�Q��x�H��Q�����|�ï��O���)�җ��M�ѝ%8\׏W���[�&s3q��웛Bl��Ko���ۆb���|w<��ClYI����4��bos&���x_t�aGcT(�٦υ��������vr�Iꚸu�\������On��i�]�w~d%x�)�r4.Q䣳uT\��1<O�1�l����e%4�؄��yO*uq|�|aA��UTj6Yq�aHĳ�9�}́��̦&�gD���w�bƶs��ntj `�&�q�����v�2�^	�'�2Vz侐�h�����O~�J�@ˏ`�3�v������ǠgЮ�9ª�ͅn\ko�ufl�J�q�ܔ��KC�;�5��C�S�
E�;s��B����A�n� -9-�L�#�Q���d��!&���������E}�޿e�0ޅ;�*-ԏ�/WoR=�>:с�^Wy��p���G���^��FI�'���X�!�o��D.x����c�#�7"Ұ�qa���H8������a'9*���7&+.6;�JGo�Z��0R�ל��K}��y��}h�Y�B�W��;���_���4䤻���U�b���E������p�!,P�T
U�Ltm�D}ԙb�s�mq�E ����@�l�'j:��������%���MYᗶ�6��+���k����e�@��7r���(>>��czs�Q�E��-�0s2Qd��L'~�M��i*�D�Z��d�k�jtfg�$�H7hWW�c���	_s��s(��������L������z R�[���.�FLw̾��7�{6긼��u���mί�uMQ��&0�Z�%}�X����
���Kt�`*w��/�i���8bt� ��s���+�p�Js=����Kry:��*���|�(� ܎�rZf�|yg)�>�*�}j����Cw�_m�C���Ӗ�$
����w�&�kM䆣��3�|����%tx	�\��y��y��J���.�m�e�ww��{Y�'L.OK��H(�Ǽ�����`rzظO�?x`�pt��/nS>C�.:·�9���J���p�Y�u�ī�Ӎ��O�p �ɍ� =�����~�i���G\���s�\u�� #-x�BW<Oi�=�b躳6�g%t9ș�����<�������>��>�@8b� u`r��?��
��%B�b~.�����w�}"��s�Ri1o<��I�:��v�sq6wZSZs�h7"e=޾4K$
gBpzDy�+�Q��sC�� W&D�3��ɘ�����9Q�國�#J�h�y����iH�K2�b)��5:��go	Z�	}͙7�������	�O,����5�����P4~�PH���Y:Z�ɩ.��Ȣi���L��y�=�A�Ʌ�{<@K����S��{۰���r�ɕ��Kl�NC=�WJ��Y>?�5�l��9J�ۤъ`e"�p-�r���Ɓ�b����y�xG�'���l�r��
�8���9L]� aՀ�a�����X��7��A�Y.D*��&���<?��X�o����7���[��cyY
~����R�z�(1w����4�i�����l{�ٵvW�$&��רϲ?�$��/gq|mޑ���O�~�ԗ�G@��*-�L�CK)�_���y�X|͙~��'�E�w�]�l����t�0�܆jB��&���uang��L��k%r1:P�����s䀤����
gb҂.�4P~r����-��w��F�(�Jb�-iBQ��[R�zp�+�v��c�L��I�f��q�n�\��X�p��*�F$�nЧ6�t/�Ժ�2<��|�1�ey������G�5�k�m/h���<]" �	�l��ni�BI�kS���^�h�T�<ômP}э��2�FJZ��h۔ԥ�8H�δJ3!9�	��z+?J�iw_�����8kw^n���7�c��'���v �	$��2�	�*1څ:-�GF�Pb_\����ǩ���/�]�/�v�Dn��P������mk�cΛQDԳ�OC����Ŧ!�G��U��ӝ�n�@t�!���-�~��)017�	Z�S4�Ϩ�P����3�=�}��\q�@�5Ʋr�go:i�g,�*/���}�7Gۄ�� 0���yPj��\1o8-���������x���U�x�Rټ0%���U�N�6�7�z�$4bP��*9����E���Y�".����\����J0'�3��N�C1�"��.�r\���͋2HyDGJ|?w�.�8=�W�<���~P]�,�D̴7L�����
��~�yB0Ljc�N�$��1���:������J�@��,�������{����/e.r�ԟ�+9?�[	ZrWl�w�ʂ�#Z�u�J�V)}}_ �JyG�>R�5C'��8�K��T�p<9}��?�q9�;j2qp<���w����5)m.�"RsvM��T����Qm���R>ZJ9/���w�]�}��-Β�
I}]���%M@�����=�`��:H�Nn��8��$r7�T D��\8�"ux��&���\��aNZ�#E���yHY�H�P�رL.�"�Nr��}nl�`);���\����:��3��8L��G�p��( �,v�U
���}�N��Q�c�a ��T(`U&¦J�sZ1h��:�v����p��[�2?�R+haWH���q�n�}T�%�6N�*NN���>�cL�C��6
v>�e�?�4A��E	��*h�2	N֖	ТZ�C��X�v=�,�H�vAk��oT.�I��Qm>��lؔq~I�r�o�G��	�^hCD-7�U��6��<��R�T�N	��(�]�:�px@��¤�Ĩ&FM��0���iA�u I�N$Z{�A�	%,�D4ybM̪T8���(x�ZtZ�ه�Z�c�t�ž���N+�mb	�h��
X-r0�)��G���6���-�6�Dk�8`�0#a٤�i� n�ذM��8��čaB��I���M��2>	עJƨ n>F�0�3�H ��:�\��ه��uӂ\֤�s��%x���) �,�:`]�4<��i�u p�aM�Lؕ� 9���8�:& K��	Z�3���������l��5���a�%/��/i�n�����dy� f]�%��m}H1��͑`��(O�H5�bc\$n�B!�����<M�a"�(*��U̡&u��)�V1rJ��*�F��m�8@�,I�X�xk?�����C��=�>7�^W(����,�ЁDKt���J���P�ǟ�E4.�ގd�/�@ G�Q
$-��@-�Q�;E2�u��6�\�yd����Ѥ�@5�S1�*�J��;��N�&e6�zu.��9�H�u}>��-�a�i�N$�N�&�{��F�9Ы��s�&h኎�VsI IRª�!�֍D{�,�B�m	:��`T[8����iy��!�|3Zk2�=���t:EF
)�"1QF��/��'��F�m:�3������-�㴐P�)Rst��	�3�j6�Q��������x���s��1Z]\���f��b�J��F+Ϫ��䦅V���ɶf��m6X� -,f3f��
Z��7�q�.T�b��8b��<)g����1��@;���@���J��^�VS�,��lv���&W<��'Pc�I��.D�@M.��C��.�!���%����a����ۜ䂖v��*���9�C��\�X�R�y*3�wK��7N;��c9�6'+����~���?{zG�ݫ��x��-7Hqa�s����+5Z��5����`����LFa^���g#��Ft���b|�)�E(�K���l�J����p�{^���HOBA^*��T��9�S��:{�a6����&���N��=g���k�C�i�����,,����P)]���U����hDG�fK�őZr��˰�&&�ɵYg�
��,���<���7�i���.�UyX��qZ��\�hA���:���Q���Z�v��R�XR�1�	v�u&-��dEO��M��0�䂶�4kV#)^9N�����	��ڡG[�����\Ю]U�UK16f��� Lf��EC� �{�b��Kb��rī����@�?��]�@�É�Q��q�l��]�X�	ڭʱvU	̝C@g?���ĐR�F�}F���A䂶�2[֗#%^[K��h -:�@����!����~�r֔��;gGc�)�ňJ�F�=F3��-�Q��rA��,[6�#3Ykk}�S1��#��6�80:�AB.h7�+�Ƶe����l��ܥ�7�6t�����`���UІ�zL�n�X�L��7ao��C��Y��uZLuDA�y}ԍ�@m3,c�	OH�Վ��5J��tqF�<<��P]j��FlE�����Z��Z1�H��k�i�j�`5'RsU9���V`@�C�@KZ�k���GC'����@�ӎZ��B���-����R3l#z8��w�v�Э�`XOZ�q�޸q�����x����&����n���P\�����k�i㊢knؘKHr����U"�*Um��*}k����J��~G���}�%}��>�I!�HBL�|���R�sl<`<fƀ2#E��!�u�:�������ބ��n2��&�<�9�'��<+�YX��X;U�l5�����`���l��"L~��j��b�_��%O�L~��
TS��Lʶ��fcNQ�%Nډ�\F� #Р"4,<w\�ge�B��_+�{���h�k&�$�EM��DP�1tO�֝��7���ӑ�>"}�����z�	>%mw%:Ӯ����1a񶐖�Ǥ�����"q�VZ�o�����?���K�wY]��MI�71�͝�m"-EڻW���s{&#}� �nI+��f� ;p$�4��0�ד�qvi��24˄�DC��Y.e����G˰��`����`��@_O����"@X��;��ش\<�SP���Xy���U�����`��rJO�ǹ�-��s�u���Ht��\��2
�G;����֝6�\�j^ ��x�y��f�&�nO_��\����a�;D�$,���2�Ie�)��d��+p_��Q*��/@��DQ���^n�\X��iy�=e4�%��Exֶ�H{~H���
��:��+|�۲"�X|.%��KDQ�^-Ü��W�;��I������D�A��'���tk�i�V,:�RڅWѠڤf�R�P�:��|��Lb����0�5��)��v<����-J�'S��p��`{����F���	��&�5���H��ә��`�26�+����>x� [zb�c��*��J�O%Y��XhT��-�T媕Hɇ�=�n�a�X�Vچh�~�nbQ�-p,N8i��=��2ʒ�c��Hk��T���¦���F�.�N�7��a���u�8T�ohV׫(����Z��?��&G��EXЕgZ.+�7U��AQ�+�n\ƕ�w����5��,^�u�E�H;v�,޿v������d��β]�*
u4:h4�Z���>�+-,��",4�c�U
_��#j` ��,ȑ6Y�a����F鈢6�3��̆���kZ��C��0��6��`x�d����Q�����訤=3�cs��K���E']YQI۟�cX(a���`�����z���vx�c��6��d�8��Ǉ��#�c��9�[��6�qD%m�J�$�@?3*i�ǩ��I�B?3%mٔ�m,N*iOU�8%mR���ٷ��qd��Z�i�MI��v��'Eچ�01��f����X�ӕ�'z�H�� '5F����"�E�$�a{"W�"z�#�#���d�p<X��;-�����._�*]\�k펢"O0���4v�u��q�Vơ1	�F���:��/eZ��(*�8\(8�3w�NRw9�3�������*�"�M,J������3��%!��2���S���ƭH��ދ	�W3����d:ȭ�ؕ+�v���	��4I��n&��i�)���>	S�06��s��,@b�\(<�L��8\A��Me}r O�;f��Mg�$P
��  wIDATű��=	����=+'U{�*!���H�?�l'��?��@�)�4�7��A{]�%IxGU7�A��'�t��il���Ƃ۳$��Ͱ��Ӽ쵏9v� �m
���E+�т +R�'p�z��iCQ@֭�vhE4FVf�q����.���B\6-�v�E���?f�9�����%�8�E<Q�G�р�^��:�W)�l��65f�C��Ħ�����s_��5� �&9��&��/2ߧ��ڎ={�߮���&G���|v���i�oA�'��;���5͹w�%�]�1�q���-F<��c�Q��j��6�8j�Mt�ـ��n�*�� ۴(���q,��2o#'����,b����IXh��i'�t w8F�h0��?����4�N\�C�ݍmGT��<�F�4�b�#�ЮI��0����*^,�fT�;�Sǂ�s�>'7E�6']���m3�5�^��h�a�y�CM?�"�"@��;m:%))�{�8|��'RR���6])����i��?������@iA�C��MM�ΗR�C��^�**.T�/g�ͽ{����>L���������{�(Ce�����D�u�Q�C��^�W8W~�{_LG&��Hj[���s    IEND�B`�PK   �}�V�Uˮ�# s5 /   images/fbb65e9c-f417-460c-abe8-d9c00fd6ec79.png��S0��Cq�n�����q�www
�e�w���ݽ���s��s��{�?���S&O2+��L�ʓI���
" EFZB���Bv]����tQ����$<�� ���U��?�X�cv�u�X�<7v�n��@�� E ��/�0RPy��b;��:�T}�npd\l��d#��I˧0��	�*�4�EV�u9��
���t ��˃�/q�Oul����S1X������0���1���z>�n�������/�:0���n���/q�y�D_����L��_�����dS�R;���Q�i�+v���ӿZ���g*[��X����l��n���������_��b�������/������V�t|�]h-���D��y��U9��#��v���0�8�j��~n�w=~�?�ܷ�[��A8����g	�n��g��o��^�~{�i̊�^u�E�~Z��'�唴��.|���o��By������3*�H� �lߙ��1�tM��w���N�e��� ���a-��.���i�[��7a߽T�����d�X�'7RC�ۚ���۷d,�ss�w�s��g�R�oo����965�Jbˌ|�G�υ�J~��=&�o�F����N�wrC]pb�*��<�}G� 	���� =�Z�L.�9�.�/A�����I��	w�]/M��I�7���~�/|Q�~�&�a�?l��Ţ=S�15�*��	��1���b�*ʰ��1Ȓ.<��C`a���_�X<1r�i�6q�]��u��niq�Ys��o��̅�~z�@Á(�/.��k��^�]���Μ��k��˶%g���ē�(u�Vhdѫ(*Om��@���Q�S�6P�ڹ�d�Ӷ��s,��_���s0Ԩ羌���Q�5��af�$�s��� ��N-@��[٩�T�e�J��r�����N֋�`�6�%�\+Uw��Z�U��S����i���7��Gs�D��('��V��7��c׌>�_��ܫB>��{���nE�u:oZ)-���wF^6�8$�O������?����~�˭sO�ʷ|7P��{��1f�r�q�'�<�ߡ�Q��6�:$Ⱦ�w	������ �˵�L�\�����1�s�w�w΅�l�b��x��sZ?��כ�U�p�s�?��e(�����k�_���^Ƨ]�+���I\�Q}��~3�;S�^0g�/�u��c���ͥ�]6h�4�Ӳ�}e[a���YuX����&��L����u�L�c2� N?2� �}�D�<�>!(�L����^,G��XjM;�|8�vl�xrX=���2��p��Ѐ �n�2$Wm�g劫\RY�Pu�=㣹���>�G��MD/�UA���"+�t8zg���ʾ�MR��+(3v�����F*-����Y�/��w� �Ζ��N�Ӝ�T�Q^(\H
"Y��-кv��W��~IT�Om@�D�aEZ�P�fgfV��6�Z-'�A��K���K�Z�	����<�yߔ��։��-�y0�pS�Z--
���S#�88OdA2�!�"vA�������2$vQ[E�D�@��!�_�'�k�G/d���z7�1D�s|W��2�x����*l��"�Ě�1z�����9b�����?V^lF�=ųm$�[�������vP?�Ѝ��^��4�+T/Ԫw�Y�A"��^�ʚ	�]f�ꭋ�3G(4�^;�����zH�T5��԰Ms��~�t����͹$�dr��C'`(�.<�uͶ�������cN#f��}�X�đWDу�t�f���r�������d�IG桉���4�'����=عcI@��~�z͘�uQ�l)�r_z�"��S����tHx�7T5[f��3��5c�w8Uw߻�=�s�p'���Ɉy�DsH���;@� '	!�<�-��Ep����P���~;�p~L��[�V���ư���X /`ML1z?<�RC媓k#�(�==r�)'��9pZ�L�<��ġy����Po<5�=$,��,x�
	���-�=�lj������dx��{�Fntwl�r��z�;y�f]>f;;�SGD���l�A���03�؍E�9HG�P.�I��a��|Ľ��t#I1*�w���f��KW�i�8���n�k�������x�|l�c`#t��F*1rj�<��U��uL.�e<\�a`��1 rn���.Z ����:�eX1�tgEӛ��`a���`3��g܍$�H�0.��!��e�#��3�����b7������9(�'��\��m�%y�)���Í���oŢ[��(A�*4�ό��mA����v��^v-ͱ>jk����;�_�6v/��GA[N�p���).�j�2+�r����C�cߙث�>2QN���`�j��m�0�!�B�e~��~��\�������ֈ�����=�9R���A�����U�0�լ�c�B@Co�>,�@�wc[�\[�TN+�au�}�5N,��.��Ϣ�2mD�J��O8*0�f�RL����u����N�a�^d�Z�y�o{[�])�8Jc+6)��@�:p=�?�����\1ZS�fƱ�F��d�UP8�l���fB#V*�~�.(�B7�v��6�����7F\4;v��͕�Dh� �� �uHf�=52��v*�5�os����������W�Bc��4���:D��£[ƍ��Q���̒��%�8%읊1���;)��^��~yC>��B($��;�aᇩ+���n�{7�X4./P"�ѧ�
4yN�V��ɬYO���p�	�� ���ۮ������*��*�f	b��<gv��v�x},I�����l|�ɴx���i�<|l��}�'�,H�!)�]w�
�9�1��b�~�y��ԵN/�]UC��i�S��~S���.%+j�����gFd����LUrmJ+(��[����qt���->8��r���1)��EߚM)�u���CI9C� PMA^�R8��#3^�7F_.�|nq���tmqʵq˰[�z5�t Pp)��"y��D#bu��9�E��ދ�+�x���v��9հ�����1i��%�+�t�Р��gq��̢3���H�.����`��2�B��/�۷���v=�A��+TX���������[�g�чu�F	��9��^j�,�D��T��~��:����[z#H֚/Q�)���C���W�"�4Q6`K�mOH�����O3�����޶�Ɩ,�I�P?`����0����U�F.ql;��U��7KNɇ8���\�)h 3_��ӆ��[�i`����Y��6� E{�Z��b7榬�ҶY����_��j1�����%E���P�KL�X$]�ٍ��Q���}���&���6�^�5���@����=i4�Y�{���hq�3��3�%�W�X�����i����?$o��O)���wc�	��vk�(e�cy�|���h�EWĢ �����(-�T�Ҧr��?+9���\��>����W~�3��~\�:�#<ƅ�\)L��3d6o��~*�Jk��*��cGs�y���?��1 	/4ޖr�`\��u5YD�tj1P凧��������I�YW�f����
*�箆ǯ���(���bp�z" ��������"=�»�L.oȝ#y�@`�xkax(���h����� \����q�B�k���nR�uTi|k M|�Z�� 8Nrތ�AAԦ�{1b�Y�G�O``BTq�������k��ҚeLW5<�_�DI���<~8z�+㭟q?��蘠���ǜ��*uɼNoU�����Ҵ��J/]�R(mXn��v�	�P�%Q�5�s��Ԛ�+Z׷��xd��]O5T'4�)/��.�/|�u,G{|�Y��e��f�XDP���þ��\U}%CtWla��՘�F��+����,T���{�pbZ�)k9u���T�/�\�x}]K�8��?)��k6���
�1��B�����斧N�
PY�9
@��]t^k�i��2r��6G$��wݎ�\-�M��>m7-�w 	A�cGw���U�b�:��Uӥ��#�h$�q�#܋�w��@Ӎθ�A	&�G�f���a�4Os30P_L+"v؂����!�|��CL|��.��%��XF/ �E�f�ϒ���y���`v�%
��±槿��D��W���7�-7J���|��ѳXL /������L-���'���U��w����)���"��5�/����N�����0��ݯc͇2c�FB�������"sh�B� �`w�V(^]��^�1A�^*�L��kQ%z���zLDd<L�&����E�op��57���M\;�4��J6�)QWRpD�-�ǃV�V��F�C�����&���N�C R�OF:>��/��*�V��R#��CҞ���!�n��n֏CD"����S�����q�B��s�_U�Mq/%���3۠�L���I����闩v%�N�����s��I^��]�"�(6WGc���<�9R��}�	 O�f5�G������ΥY������8��ϪQ9O��P�<��)#\��u�u�]qn�*��6�lBh֠�$oAS��*�Vפ^����i&�����k��^Dn�h��LeVl஦d�R�H�'!�QN�t���R��O5|y��� >�s���i�cLJH��V�f��,�����OC�� RC��OHF�r��q�$�H$a[��.��r����d⧃Q�yh��{f��
��s��M�����v���=���n߹S���`m�(���#����o;���&��Vb��P� /��J��iŎշ�ĭ�ƃSPD^���f)�S���Ė8g�M�GJ+Wv n��CNr��m��.ʜV�n�4��S[����Sn��SՎ!��:�J"X���bX\��{^c��
�^=��.��A�)�q�#�1��I��D
4��nC�į�	���>gV�pS�D�e�'��|DۣW,�`R�~'f��Yƺ��f��\5J�f�d�H���E��`���!J���5`���$:	a��K�_-��v�� k�{O+���Y�W��C5��o�I�SU�n��ߌ{�qpn���&�,�����+ �:4�~�n�p�hT�r i0ph�R��%l�<Ct� ~2�����:��O�[|��o�!q$X�E�Sz6ו�bˠ�2 'JD׫۠9��uv����p�d�Z���@�]�/dLd��o0+0�]QWx�㭈���H�<0�۬��v�Se�ig�K��{����/��Ο�،I01�k��4toO�� 3'op��Q������}I�"=�.-3s��('(��./d^v8m'#�%:����ޖ�z*u��q�b���oI�p�����n�'����Y2q�⫅ߍ_q�'qeƌ�P�����'�R�(R�撢*'14aS��$��t}�Y\]��[Zdz�E�	�9��H��hg��$��	���;Uc��j"��"��F���}\7T4�K���l����١r�m%*j��$Oc��Ì����Wy�����qػ6S2��m��g�a�Z�ࣔ�U2J�,-��"���������I/$� �i�U�/VK�eVu�CT��!	t����;;.I�`�]���bm��gqj��(ڷ�p&��]�4�Xd����
��@��{sqs�abȨ����-�{�D����k�e�6ÿŅ�iɏ)���T������b������^F���EڨnM����d�3��F�%�y��BH���Vo����'��bv^t�\ǹ����j�t9y���D��&h�ݸ�����E��U������q�����&K<�X��j����#�u�8��\�58:����I�\�O�Lv+��_ �v���~��cE��Gr5���I9�6{3��?땧Y�6E�3��+,�3QI��1p��u�[;�y��dʓyլ��|�
!0ib�b�,7�r�c�$�u=�onw,v���u:��DbgsI�|���f1�DT���Gdp%?ӷ���<Ӷ�@���޾�M���ư��ZV%�4b����N%��8l��+؂����-~U��}�R����=�H�tpF>�-��x���n�ۮ��I���TKy"޹����M������+k%k�zxX�S�?ԥp+|���]���{�P�ݟK(���ך:�����_��c��IfC]�*�]ah��X[|���z��OL輻�Qk�i�-xOR����h�_�� �r��F	gF���
8ڶ���2�,<R}�����,�W|�N�x�T�����v|�;@+��&8b �)D����Vy��-���#i�ex%_|����G��q��w�b�I�p湽�G���v"��џ{�|f����YY�%���r���U�5�ů�0L���(pȍ3�����=S( ��Q�m�N?�h&?�kL¯�X�R�dQ�SPHȒ�w��1X���qpe_���iyJb�["-�6w՜�IP��劀�ls�Tڅ㚕�q|s��fyo4s��(Τu�2Qb�q�� �t\����j4ӞY�s��H����d6��z�9���ߗ:���K�[s��:kn��NZ���7�r��%�j�$dU�ԕ_�)[\�*N�O����]�?sh���&S��U%]�ڣ��i�:=�T�D���S*E0t��=	0�KҘU��?�v�/��W ���`��h�D��zD*�$�^H������\e�;r�3���ԅ��� �ᮄ����B̧���v��$ �TQ��	.,`!�`�QZjA}9��'0����E����ǫ����Ǩw��$rZ��)�AP�fPB{�^��h3�ƽ��i!�.�����(K�tH�;?	,L���t����\��
��x���~�e��|����]з�qGg�4F�E��hv�w��=P�2�͏��D���Vx�o2�?�RE7��]ڪ)�Hl��6`8G�����\�\����)��S��#����tך�tcpް�J\�DϬ��>b� �իϢuQ\`e|���"��(��� l�C�1�wbf�F<�>�:���\�C��@��ŬP��A�\4��������U�:Or˷'K����r�v*��%	���8�BN��_����+_Sřa++���e	��-���	�{9m�ʰ|I&���s4�O3�C㻲��.���\V���������7��r~�η>_�L�:X��� ���=�7��d��2�S�'i�F �d��`)*(^��!��1��/�UG�8<��CZ*�ag���f��;G��C.��H5Rh�$�e+j%�j�o�¼O��L�L���p'dQ�a`9�^:;�V��iLA-�[��j8n�E\�WC��q�����5������B����I�r�/>��	)Yx!^#+W��5m������g|��GT"�Fm+B�����L�+�}=!���eq��lÈ-�N`R]��<��7���څl*��4;�U^
e誟�w��sq��,-�X[Sxa[��hD�=���2�Eel-��j�����%�ߣI%��U���� ��?�}n��3����QX�-Z�\�ȍ
�����;G�m�*ic�T �ڞ�y�����q5����b����ey��ן��/Y]��~�p�<���[S1̂�Tՠ��֐hZ���_Q�.�PQ�Q �.Oj�	|� ��Q��+kbÄ�2]��W�����N�34�������2�?B���!��ƕ6�@dNV���X= ]���״&X��a����2��L��k.�<]ߗ�z��Y�>3Nv�|X�3�W��#��f�T�B��%�q���b��p�-W��ȍX��1�e6�p5��̯�o��mؕ�Z��N�+5{�6��k+U�{�����ȯ�n�����K{N�ns׶�Q�w��e����,�Ƕ9X�h��D{nL�B��V2�c�}l�0�����_U�0Y{IJ*�|�nʤ�����`ia��R9Hs^J�$��x ��D�jz~F�,F�I���b��d�T�P�3��^���-��A�W�[r�j�C�ћgĶw�V�^Z�L����;V��<6G��Q�Cr�?��6���,�1�-F��*�\�l&ö��-?3�t� �!�s���n�-��n"�14}B�7h߂�eS��� 3�&�{k<���t��	����f=8F0poF
<����G�$%7[݊D/2ݻX��esS�����oj������?�ʮ:PV�LW���1�I����>k�N*BV�td����>mN�:d����-�?���l�3$V���s� ^`���
X��!���c���l��w�����5[5�������|�mWK�8kxJF*�F��yƸa8�S��$���*��-��&;Z9���ޗ�OJ_`6����eԚݓL��l.��¿k[�j���l[H��ʆ�3켻y�'(�e(�� �1��P�u�]W���+�c` /KP�+T㡣@�dF�#�2�G9]�|x��&"#gy�JȆd���;ע+�	n �[�q��|=��L6x�'י�2��jx���V�Ys�q���l�`N_>xX����;tU*�̷�,�������G#�*�oJ�T�ׂ���SȚEC�?_&%�b�1n�<:L\=+�_Z�� []�[�̶�~�s�>|BC�A_�Z���Xu/9_�����k'���Z" J�g���rZ���N��Q
��4j�L��8|5Ke:�s��pT�����B�ʂ�%U�lS"�n��L큷҉�)A�b���h�\�	��,�X��7�%���1Li�4c�w��X	Jp�͔�.�U�9���EE5�s�ţH��6�y�\�xE�VVU�t�(�w��b�S�vZ�>0 I%q
~�4h�i��7Y�ғR	I�YC��w�b�e����9�T�,�S��I_�A`���TGPM
!m$]�u�n��ȰDg�ݦm�B!����П�Bh�0�w>�����P�!�����u�Y׽��]�f��gف<�7�-̀v�N��%���}f3b�5~TS�R����I}���,��"*����!^��X{�{��H��t��̆Ne�Z¥�`�ۼ+0a�Y1@��y]ͦ7���ƾ/�g���v��=����X-��_>nO(�4%�.cОc;�؏f9�e_ ��;�{�8N������H@�$�[D��|W5	�a��ݭ�zw�X�b�`g�9����:N�ᠠZۼv]�������K��m��_��Ɖ#��)u�RGO��db/ؼKF2Th�)7P��'#���%������|A�)/>Um�m�|.H�Nr�vfwl���^�k����Z]�-B�R.,�fa��졦W�ƻ�&�(f��l��t�m�P�ua�n��:5M���� ©)��DUTP��?��K�������6���GV���K�K0M�[��&�j�JD����Yl���R�uk��J{�[0}���SH�]KjPшP��ޏw��@[�0���YF'K���E4�2�f3���H1X��v�f۝��&����Ǉ ����v���b��F�r�-b۰K����w!B����Oj�,�swǳ=�;�����*F���I����vc)<+�i�^��փ;���fO?��Q���HE���1�,�0��`�+�U���K��b4�Ie&W�/����[��+L6O�� ��
�g���[H,�ˣ1��1����Ck��������O�·D�f=�Z�SL�$��dNr"�A�V�N���bs�ԄX����99V���c~EX�ů��+����vX	ki��͸��`��u����
��<$<�Y���r���%�T<�c�`
�Sӎ�<a2� ����u����&���?�F��W�-�\v�ʻW�G�}.�d��9� ��T�W�æV�Qg��^i�̚���0�QEKbz:�L+����.���"Ϩc�yS�z���b��Rՙ�%ݏ/�2!�]���`�xcZ*��H���l񨹹�w�?�o�u`^�U���4ݙ\���)gG�^9W��Ķt���laEM�������
V7*B�JKq�99���Eq���j�R�X�IIw��%��
3��B��E�;�CzԼ�%2�V�$z#�6V9;��B���-[չ�8�r���cnC�Q��l��ºG�DQ��\-J�TeV�$���h�!;���w�DD��i�?@x��\��G��l�{�I�ݞ(���8��L#��Z;`';"�&��[��V���}//���ճ�Ņ:�|Dу��"CF%L�t_���;��Ŗ�[h�l��/�)���-����F���7��{=l�{�J ���Z81�pk_��v�{�tq�ZY'}��-��U�@�����+;��Q���0�P=f�N��� \|4���g�vl�=��x)Y�4%�B�'�����(�۷]k�����x��j��:��3�Y쫶�=Q>/c'�Ό��CM�j�����V�����P�9(,y
��~���W���fIs�"������F����K����,JDF�u)�s�z�f������~_۰�y8�6��i>����dͽ�� ��hR�Z+8�P��"b}��θ�=�'nt�.LBB�T]���b%�V������s�#�]6wm�̙�
��2c��/ԗ0���^�B�(�>�U]eXҹ��������j��;��;�B&ٍ(w �J�_�A@5��Δ�<�2����huҝh�ɖx��Y��\�U�^�zRt$��.����]��Gw�Թ�v�u�-�"1����>YL�Rt4���˫���/,*�n6)����I�/OT/9>=���ڈ.�Ėh�����M.2ma2q^Vs�`2��|'��5�Q�O��#��q�z����??�M3�ʄG�R�F���"��8�O����o9����I&ŜSR�Gˈ1�FE�r0{��;[���[o�5���l(��d;#�X'��	���������swJ�ز��<;�ϋ���l�Q�C�"�������yՊ{���$�M.��2sR�@���k6������Da��k��H��d�m�S����ϧi�~�x׽�<.f8�l��Ӈ?��۫�����&7����9)��T��~D=)	GP+]��Op��e��+=6,��u���#�]j:�cC��_���(}������2���	��Gy�z{7�p�s�Y��������?N{�t ��C;�L�~l��`ٞ�ƬIg�v����{��urqJyuy�+�)PYFI�����e� ���-�֧��~l�U%Y�ffip��"}�]�U�O��J��S��q��àr"��Y;���Bx{�]S��t钷�4���9o���}aE�Q�g;�����\��]<��c�^^�B±�W&=�A/ڛ4^�l�;���<He&1�3�<��Y+S��h%�_���(P�ѠeQ���+�X&��k�Z�q�G�5.��or�q0��>���*�B�4όH�7c��8��in-����U.�^�f�>�r��jGc����J�XF)�E�tw������<x|N�g=}������~w�f-@x�l̍}B�+�L(��Z=�������'��V� �;�-��ޱӣ�aГQ2ۏ٢�gG��q�^��A�r{3)�)�9�sȷ��9WpE�l�L����1�⅃$�����P��i�S�� `�~��S �~�.Ɍ��i�U�-��7����
�����o���wsG�� �K_��ڏ� �<
�k'�M�2��(��+&�;�sh�^^x�܍W'�����k���/���Ef�'� ��6��Ag�|���L����VA�+�KR*�a�N��.�G��Bo���D��i�>x��v���jSd�[���lj�fc��n��X6L�P�6X���/�u�T�н�/�i��MC'��Br��������g|i�t�E1�x�Y���֛����� 9�x^,r 
rj�vTc���K����.H�$�G�Fu+�,x�;�TT�T����bĤdf��>���԰�n�pQ�X��|�:ɤ֩ǲ>+JԢ��d7��CFBv����&�`bu3��<�$�KP?�{W �"�/���@$A�h=��Er�@��#v&0Ԟ�`k��A��&g�
�eڜ#����l���*�]s�a�EXkr�bֶ}x7~4ؖU��;)P?�$�~�՚W�غjX��EM�0a%R,6=U�="��+U~��Ђ���U�.�9�|�C�`+�1�Pͱ��jw����4���x���Dŀ#_�o�*y��r���[�^,!�}��%"�J.�t�U2n�a�VIJ>O��eN�eF�m��W�p��c��{�dl�
�L���+Z��t��[ͽ��&_���B�"��$��K�|�^����w}0���2+Ό�B#qS�<��(\���1%�c��`+%�~�1�i��#Y��f12��X����w���`
ߣ㦦�_t|�+�:��mBW+�Q�j�_�z�=\�U0`�����V2BY�H 4|mK(��V�>�2�"�6=������_A�ϗ�p� �ߥQF?�,)�Z�y}��������Q�g��6�>|�[����Z��c�~���ܮ�^�+l��t{����1�J�<�Smd��EW.dP����`|��V��&Y��9���s�ݪ��[=�Κ-ƀ�Ӎ�TŔ���TB��V#q�p6'�a��7����~	y�/�����]9l��ܰj*�F�ڠ��t}��&C4�%t��/FlJE��m�ov�!��35�[�g�O(f��P��d�J��M�f�Q!s��շ-V$<p�Đ�^����N�Cn}i���S��{��۸B�X�㏇Cy�iǄ�9�0'�)īg1'�9�s��>v��.��B�Үh
�/3��Ӂ�ƞ��t��I�Q�5^�� h�w�V��r�dq�X��Wa��˶�F]��>4�4Ո)*�6�
��l��'�;��`�2�6ld�*�]dR?�^�YA��J���%p7�3��k�n�Z��4�rr���^��|��
�V��k@iWqW"~��2c�+]yl�`�����M�aDce!����B|gF 3��1��D��LS�p3ll�Y�XX����d"� Cvq���'] q�!�K(3�����w�mp�m�ĬPc���=+_�`�q��+B�q#�d��dJ�ޒ��0�Y�����cu��8��B z�ɰ=~��� �a�f�+.�m�h�weԀk�F��?�;J��e�_����X�����Sg8Dp}<�]n:jOYR�?^s�����>BZ�^����:�$�,	<�]�c�V��|X�j��'��ŬP	��j�Mp6�?\T��GbČ�R��=c�@�~?��	��� �JIP=��R#�4��V��j��v���w�-4�[l��;�$���#C��9��5P�_�d����"��}y���t9�R�-q����t�tx:dڶ��=�~�Y��tD�v�G����$8;Tc�I��L~!H�@�(Ïys,��	�)���Y�z������5�D����3�[�=���M -�V���@wy0 �o�y[q�#1�ҡ������Wɸa'�&EZ�E?+����3_�yc
���t<ߝ�%"i�N�GNJ���2W����]T[k���N���C�H͜z�3����DT�LG�^��S��������%5Ԧ��P3Ґ%'Lj"��J�M�xe�Y
�zO�4�Liv���:DO��L�j��8y����	�l���<�����i��=yфV�s�(��.ꂤ�6��G ÷�n�k�rW�6��9��b�c�L�~��L�2 Ǒ�_$��Y�^����NBi���jR��邚[د	���0�+L�%�vܒ��y�)��>�#�Vd��k#_��Y+w󯫯ɹf�j�q*R����q�c�^��_l0�p��O�;c1aŤh�W�ܖs�i�)|�rd^����#�V��R�#bvb�r�Iۮ$�AP�=i�BU"5A����W�
+�V�G�J�Pkm�q�\��	�*��/�_8�Q��̽�_:&F��iJ�-4C�%�eA��sv������ Ʒ8�m��`�6�0��L�}RT�'|Lvo��֪�ϭmG�?�nܨ�7���xS���m��PԊ�}�}���]�!E�=��;�B�2��WB��Ð�����R�l
�qM�Ǎ�X��R��hV��F�3����M<o���<�v�bu0^���lļ��t��}��XI�|X�l4;Vo �T��ԭ����}�[؟n7�A��c��=t�ޛ*o�}m������i��5���f(C�b���̺�`�ራ ���(� �0��vv!�  ���������m�$�h1cr���,/�ٞ7A�o�q�;a�el��j����Z�����OԾVJ8R�фHN���@����|���I��3iv=,2� ������	�Rs�ϫ�+�j.݋����e�qz����ǃ���y�{:G�!Q����D���㛌?jqJ���Q��1��q��Z,����<Άh�ZEVdX7O�;3\XNt���q�����(�ֳ�^�C�/ ��Eɣ=����.m�����	��.�[����t��r�b3X@$_����cd@[\�0&$��Q"�w���qli�bX�Qΰ+D@�ͮJ����PDe�\1ҹ��z]"#��xX�E��b���5�<א[�L 9�Z'af�%��t��x"+N��?tj_wé���r]5��]���N�9B����'0�N�u��)��/]�ƻѵ�
�wWd��n�x&�Ò"���+xΪ�q׾lV��)��&�e�@� P�X>u��� ������aT����
�i&�������8e*�x�Z1`��ma:1N�Bt�����N��!o�,_�O,�ζ���-15����8Z��-�N�`O����]��q%!O�I	���s���F�]�7ϲ��6A�����t���驖d�ڬ'.GO��Nt�k�������� (����!�%��j����A;�G]c�聞�"z���3����W�{���GaC�y��}3����]c���~K=U)���6�X;	w�,]5m�-�v{C�����|���?�r��W$��<o�û�a���i�?�\�&l��+�� ��^/Ý�-+4k���"v���/?�H�p�����
���5	�J����ڳzv]W]n����ӯ�8���8t�#r!)
����1��%S�y�ή���&e�����mSUq������1KS���޺�f�\�C�O�#�/k�n� �Zwz3����3p�.���]��Α劫�!�J��<�f����
��>KY�|3-���%�dWנ
U��t�[�z���r�Ŏ���� �d����	�]����<
�+Ȥ���M��7�c��9�1ʘ*���,
�����@R�Z����QX�p��YW�5��̃�פ�����ic��Z6a}�nn�=��a��	/P�=��������x2��~�1��D���"n���J֛�9X��.��5Ѐ�������k�KhĴ=��zB����r��DT=X���`�b��'l�;���2ɞ6�O'�������o}�e	uF���7rᯪ����Y�+j��ᙤ;�a���!x�0}R_�G�d�L��kaRkL{b���{���߸��F�_��8Z4���&��m��~@7#��C�T�b�����Xh��v� 6��R8��c��]Y��UX�tSbj���� �=�3�������tN�5ǲ��R[5��M-,�	���(|ppP��B-�������w��2�S���W}��Î�絤-<}�����m	�(�4�M�:>^��`�)a�,��;��@���(���������(�8�@ d�׆�����[ϩ��ZWi!�pU���C5����<�a�{R���t�4.E�?H����-�tc�)E��hE�|����ga��h˒�aE������s�g���k��v�Ac��O�.J,�tNd�����C�Gki� � Y���4�wO%���#���̇�d���%��cpCv�V`e� ���.]�@�O�d�x�d2��0�BL�͞��pc�`.����?R�����]r�4f=V@��������N�r�ۥ��,�̴��5�R��Jf��@���UU��̉P׭ߔo� ��{R6Tg!��e��;�?rS����J�P%Q���[��萊vl�YS��JYu���йT�&����U�d�c{42�����q ���~'��U�U��yH���!�#P����b���)�t��3�>I&�~�����|7����;�(�ML|�3/F�E�b�]�_7��^�|���m�?�U��G��Q�����|��
"r�g�J�s��l�t�MLELo�/ 2@Ϳe�:���zw��b���Qif ��5i{M��B߹*eP�?f~0g�t�\"�5�4}�>���ދ��m�����k%2߂�`��y�������G����V�S�����0���^O��i~qA���vhan��[�2��0���ÛW�p���%=�mro</�Y���k��u3�Q��I��6�8�������o�a�}\���\����1�X[���ǟ��c�����j��k��Y�I!�
��]�͛����{�IQ���:��x +�?�j������#�-#j/bc`,௿�������l�!��Lw�6��(��:Ǒ���3O�#K�����Z�W��l;x�0򮽴vb�(��~�BM�%��������Z��������sϼ�o퉱Xn�;_����F%�bT9�z���/kz #��4i@DcG<��ӟ5�b�������1=��t��QI!��-��M�s{kS:�lop��]TI��]��'>��k���7�����d����7�E���� aQ3�^F�5�W�1K@�,��;���QQ��DLȠ<��pR�PW�`�?7��a!z)��0Mɡ��<)df�	fh=��7���K3p�￤?I')/���^p�OW�T�Gc�`�M�)ӑqkW������L�f�`��eܹu��YOaX�XXXD����-덳ob���صk�D[:�\�a���z�~���{wY����c#���@kQ��Xk$-u�H�_#�NMI�ZF:�tf�TDV��{���
A1�|\#[�����R7B7,Q��e
��KG9���<�:���W���qJ!a<.1���@ûv�B�C�b�V���=�|/�>yuz]�>̑.��v����e��F	j�K����H'/�H����S�ȭ����trL�rQ!�G*�冺�l���]�ȣ���}�z�܋R�&�-.J���.���`c���ݍ�G� H�T��ԇܾ��4E��1	^y�ul�FX�([p�� /�yQkIfmH� iW\�@Q�L�b3��G��r��%�bn�;�O�~[j�������_Į�$�yB���Cx�ɏ!�������uXp��&�`��w.ac��W��r�:uJ��]������?x/�~io��=E]��s��ʵ7��y����+�A�;�I��q�w�$�'W�-"|�l�_����kO�n�_�%` �%�����/Zs��^�7�;/E��"
�ƛ�̓��c-�^��x�����9��i`8`eqI�۲���z�VH�,y4�Yt�͟hX�ّzf��?#�ƭ������N�fgHb����<�qg}���[}<����(H��b.`;Z�ō�z�nn0�)�Ra�p9�BU�Sm)+���Z���q'��E�b�7]�\:���]�(_\���7�MՀ��x�%��Z7O2Mqjұ�n�՝�c���9S��H�FS|+�J�6\*�?6����6g}D�n���������{������W�\��<S�Z8u�i�4���ص�������D�?��wo^�Z���p(��[��/��_İ���^��_}�;H��"׺qer]�A�oF�J��ˌ�q�ːÄQ&����S��mi�*p�#;��k�����
���l������~������$���q'�X���Z��X��P�֧��]��vҮ���.>[�t��XG(�6���^$�~�L���fʙ8R�U������n6�������[%�Q�H�1�s�>|��~<��Q߿�V���9YsK+8��|�;?�������x$QX
�t�<y?n޼��]x������+���]|�����\�~�<��a��fx��]��Et斱=��0���
.����J	�ت��)��x��"�U�o�˟����_zg^~��:�E�U��=����)�χ����7^���5D"�s�-\8��^���I�^Vd8z�8v<����wq���9,��go�ʕo���V�!��.@?�$�NZn3Қql����'�ă{������,b��E	�#0��������K������;RP;(T�|��7$��f��� �\5��9���xh9@~�֯�C�]Y ���̰Ⱦ�Y��H;�̵�ޑ݁t�e:[^b1�G
s��J�ISԜ�PHe�D��i'��Y@�8gT������,V��㽰����#�;x��-��\F��/��?�����A�kBt;>eE�F9c�'{�p�T����t���_P��	|DA�A�|��Д)i����;��@>����\l}����{�?�I�j��S�\��fӻ&�w��j�C�$��(���'ƲM̕�������+���O�?��O}�~��]��ǟ
^x���XZ^���nZ{�䱟����b���o�;�,H�|���_�>������ �E͢8��(����9��ɐI',|��*��-ӧ(&��F��o���g_�r;�7��>�Į=����:����\���J&ڎm�XR��:�r�X��&lA����F8��_�"��,�`ѐ�����	�`Ș,S!nw1;�Ru�6�%S�8�]�t�g��v��!��_4a�ݤ�2@��bU��io**�� �Ƈ���G8�0�r'ƣ�S�?��8��{���z�����s�_�
�<�#�JJ��}��ҕ�R~`�A9�;�W���$~�S����j���z��O~��W.�K���S���֏��[�v!�8l2F>fW	6 p��2|�ϨA�B�ݤ���S��8�X��>�4Vڛ����G,�0�<�!z�s�X����V��&�q��_�ꗰ�����s�sXXރ���������C\���}'�V�gn�����x��d�2�du�a��
�Ўqߞ>��Cx�}K��u|�ޢ�����^o�Nޱ��D;�w��W.Էo�F;�!`�Y�,
�����`1��W������x`�B~�l�8��t�q'���ݻwK᭔@%�I�^���tH�:h�`�+�H�`����W;Md5m�v���ȇ4�D�&B1e��H&�[["|FE�aQcߡc���x��:��2��#\�J�Wn���v?��%�nzrӊ7r�	�H�7t��7��'���y�Q4Y�-�e�Qٙ�+	"�����K��\�����i;�jt�3!c���@�Y��ֶ2���5Ӵ&ݍ�@X<�1
٦+�ej������V����RC/>ۮ�ڳ�Sy�n��xhD�+,�1W��?���𡇎�_��O��o�P_�rU&;���2l�5 O<����q��%��=�ȑ#x���;���.]��������c%8��S�p'�_�(�E���<x�aϪV�Zؽ�F��5�������� U�����oss)�ˮ]�����w_Ǿ�,���U�����!�}-�e�#s2��I<����h�7׌̤�u?l�[�**D$��Q�>�\��ږ����D��Y/Ӳ�Xuo�]�Y܋�N�@���ܯ���#i�����4�&7+Kl��k��Hm��
M6�(L(y_ŭ A��g>� >��'�g���=;��o^���/�{w��|oN���ko���p���OH4�?z��1<��������۷G��g�[�{�ř��p��&~��-��_}�����2�q[j=��BaFO}�H*�g,���0�d������%|����{_��_bi.�ڗѸ@�݃O������V��Zsha6ؐY��DY���g����U�>}����N���S�g���^�Z�F{�$��^����z�n���%�}����
�g��=�
���cx��e��U|�Ȼ����d�����Ӳ��	��t��}��q�u��（�<{��1�KF r���Oޏ��pj.Cy��w.����h �M),v�,	�q_�tη靥��D�i��Bd���#�%�!癴Y�\pvZ���m�5��fkԢ�]�*��A�e9�T�ǧW���Z�=��"]܍�^�z��w�Z-�����[��Й!bxQ H11�9��.��t'ξ�Z~�W� A�z�Q���u�^��$�Ҁ8��p�}kO�Q�-y�����8'�u�n��P�荦�HZ��/�~҈S���O��i���(������wL�Ù�IJ�s�"�.Uk9���8i�t9��R<¿�׿�?��x��}?������[7q��5���+8r���y�џ�1�]�������3���G�g�_�e�����/��Ԁ<��Ӹt7���} ]�ּ�0�e[��'�,I4c�֪��y�v"I�P��Fa���F	�0����կa�¢4Q(+�uN�;�y��v4h��\`JC�p5�֓�t�r�V:ӆQ?�=�����!�Y��/�zZ��o\s�Q1�G�nan��KX�}�q)�ä���d��`�-Ť9�;htg�Iw7������H�I��(lK;�"��)��]�*�}�'�G�y�����\�o����{��!�����1����ɓ��׿������'%�u��Y�-�!k���S���|z����~������[w��٫��?����_����#��Mم��������xfo�ˋ@9D�oc�\���x������(�n�_�/8�o��Fy��?�Vx�oܹ�r�v�&��D��^���o������ ?����>��Io\�����U$s�eb��x��m|�{�1�v#h��*#DE��^�C�!>�������H�u|��������V;A#�S��8vU��/��ެ766ЊR� �ɂ�/��,n�C�'� ����������3ܹ,����P�j~�[�x�����{����\�=u����J�ծ����ml���c�Kh�B(!�BI�� !��Bu��^ܶx{/ڕ��JZ�:�>s������58�O�؉�Ə����3�|�������5>J(�u{j����\uł�+�O@.k(͘V�m���_�&�
?9+y4
4#w#j���{-3�MZ�,���d��ʚ��ga���Fa��
�:֍�4Mh�.�9qQ�gr��f:U�A5�D����̐�x_�D]�lp��o�=���M�I���|R�T���GH��'n�'duK�#ф��h>>
�IM��2jt�$d:/E���i��e�:O	�RC'�u.����o���:j��t����]���t�' t\4��mn�C�����|�5�����O>��8q�8��)?~�npc���|�c��7���+Vp��-7߈��W�`;������ŰlÕ��a�GQ��lv�ږr�B�$c��X�RÎV]g�� J�U@qX�A�d�K�'��%[�|>�P��Z���3HDb���Be�pe�uFd�@S?rp
�����	,\��m��QX"�֧醗��^h��/�'Ų���Un4�0bճ�CD��`�.�ȥ��49
䄪�{�YvQ(��(O���h��̛��Oh�a7$�Dݚ�癲]��X�yE��*�|��I�_p���8%�09:	�����N�<���!,^�s����� �����Lbx�kW/ŭ;v��_>���&��șX���8|����Bha@2������5�"@�3֕��>��$�"�_P�-a���5X����<���	� |��,ì�/Q/�s��r[ý�Dvj���*��˛�    IDAT�j����wc޼y�w)l�q+J�<��QD�0�w E+0TP�#'p�U�d�_W4%|�q�z�]V?@�+O��g�&+0@^��u�~�
�]��ϡ����3';�ؑN� ��C d��YXߠbE�k��}�({��s��~���xE�,q�� ���<�-uͨ��GuMb�Jv�ɥ3���(��)�R�(f�()Y]�"D8@0��P�q����&g�W�-�"](�����9x|�	��I'��'.a"Ky����!ʔ��m�%~?SH8]��/��N��}�v�����O"`ң��~�yv�dsL����h�"�a�'����D�%pS@�'�'mgZsB��,I���� �V�	 �&����߅B�ĥɇ�Q�L>v-*C��x�X�^QVYDAzdKBp�sa+X�>�F0�FVr
h�(x���=�]�y�����{�~q��a�4�]��ѣG�~�3����$;
MV���b�r�b455��ӱc�p��'O�f���nAۥI<���i<�6Y���I�X܌���0�!�)b���P�O��5��L&�u^�|%�,\���s����T*�ʊO�~���)Q��WH�mh�D* 0�v�e��9�&#�]���0��;]�iN�N/*�[o�D��3a���&�GM�� ]���%���綴�gϪ��oڶ:��B���?bc�<&�=5��|�p�O^���N��jؤU)z���EYgq?�F|��@PX��P�m�ফ���5�[TgO�`�����}z�S),[�s�63������E.[@&�f�$����AXd{��#�0@���Ņ�1,Xq5N��ȹKpl�X%kƼ�A�r K= �)Ą*�Iض�o�b!��j�>� &�F�4 _�P;o>Vl�k��9#��I+��!��LL����X�b$G���X�e~�!��@N�`��p�c��3�j%�F����CmX��7l�����'q������v��f*�{�̜ҙ
�g*���&����2���=x�H2�B	�
�(a�jll�cMc �`;��Z9p�fZu���x8 A�r��4�Tױ�*m����p�,���ދNꢘBOg:;�!;E41�e�#�ÄB��y�&�d�b
V�q�u%�
n cE��#�'��M�Ia��Cӽ�DJ�(�P}:�f���"��e�
7�����y_`#�S��'MMC$�jDH��ٸj�>���=�79�Q��3��{��9�����T\�	
5�4U�5>nl)� @Ӓ2g����5����x�e���_
���7(�̍���?�Y�h�� ���i�$�������Y�X�kw���cw�� ����0�z/a��g�Τ@�WLST�������цR>���z��@8��]�n-��;��g[��ކ��)<��$�d?;���%�	��r\sWnX���y1����Oh(��JT"�`r|5uuX�f㋮��|@�ٷ�.·��]$����c<�`PǢ] Ћ�t��ɥ�B<�|�.���R�)�<!�B�ՠ\�p����e����gl�PFss3>��?��W^����o}Sd�Rh�Հr���Nbǭ;p�ny��|����/\@Y�gO�#�0���4`� Iy�p��E�,�Ű������7_��o@smJ�4?��A6�GۅN����V�2�Dr��$T���o�d��(;�I.,��Tr�.-�����,S�n��3��5�F��	�X��C|��M��T���YPEsj��!��ۏ�1R��_���E�#�h�������s��y~��~7;�+�Gz���BH��z'�Êe+��@ѵ�z�&���#��ah�(�J>�"�wz GLȡZ��/�}��a+����8��glx_I�|f_^e� ��6��/o�PC[�H��`�=}�<Ў��@�҆U �6/��� �6�`�c��9�SS�$0��h����h""�i�<*�!�⨜5��E����9�^QΧ02<���m�E�'C�}0���@G�@I�E���L�D���s`�3��cH:!����'1��FoZ;@dO'q�$��2�d��S�I��NYD�R=��/����O���(�N�p`����V�)a\��F��A?�I�P�eQQQ��P�,�#m��lUG�l1�ߥTxݣ�خ� ��Gڙ|6ç� +J6gW�2M/���l��,(�Z C�8B�d2��b�4/2t����ƳC���0$�x~񽏣�7���{.�R�s���Vzj
ǎA�X@CC
�"�����P �l.��dc(
�%*87c��m8v��8��W߄K�y���݀�c'�-�=�.��[�ێ��3�j�*��/֓<��C"�Bu%=4	� �U�^ܘ�t��b����r�v��W��L:ǔ|S`۴k�7јvT#}��r���2b�0��0M�;��5F ��=��?O����"�,�I�@>�S
MƲeK��o|���]��=�]^��s�m�y�l�v�������9���k�,(���� Zӌ��a���Yْ �ܦd2M��K�F�)f1����K��#/U�Ca�.;(�(r�L%��g���%��TVU0�JM`rb���(d��U�h��>�f�߄]��pi(�@E-y�,[���՝��a"�@�ዛb��Џ�M����H�y�d���%[Ѵ���x���-p��Js�B���Yt��bp` +V,��%�ڶ���ũ�mUV#S���p��N_J��Ơ*���6��
l_��0��+��P��'c�}3�w��yf.��
�Fη�	^y-۰d�`�:с��;�Ѣ���BVO@�.�ņFkfa��c����(�K�!y�NBh�E0E(T���K�iB�i��t�cm¶�HM�ab��?�(~U�5P�˯�H�t ^ �l�D���s���]�U"�!��8�6����	L'bS@Z�d���o�Gn[���i�@v���xA�&N���葧R�D�rپֆ��C�=a8�a��C����#CP���u���a�� 7�X��)@�b��٧:���q�G�"����|jpY�m� �@��Ե|z
~ME��qr=}M>8}��&h�	�b	�|	�D< �l��g@�t�s-�����"��Ԇ'���3@.�ocW5�kP�H|Nxmhp��7TO:��T���q��C�1�`dd��	��>b��W0(:u����5���w�E���Y,nn�;���<�뷬�=7n�5w��	�!���Y,#�J1 Y�v����}Q�~:tgϟ�5�_���7Pʗ��^�!Sp"�HCA�Ҥљ���j�D"�#A�	��Av��Xd�qyJD�LH%{\�T�Q��*a����w~����Q���¹�V0����m��6����C�C'Z�{�x7rn���cʔaK� r�4��)h�&q��2@��(�	7]����h=��K�B��4���^���X6�~� ��B	岋E��+Q����R����aHM�,�|b7��V������H�Lj�BN��x��BeXE�(�.�`��J|�ߎ��E|�ǫ��\u��"�}�Pw�)aR�P���1$Xf���b�SMc5��Z#^��?�0��a��F\J
�;?�ޤS��$,,9��櫰uq�"%�� ��b��k~�&�w���ߛ��+����s��(��_O;�_�=��@I��\FX2�eA5�5jk�c��)O@h��^�i'�O��n����f��|��'.
�a�0CXy<������*P[�@���*�h��~�TF<Q�DC3}� �J) ����0��އ��1h�̓��.#���[�A�e�U��L���x�^J�t(!OA(��8�N��2�~���j #�V�-�r�$�w�Pq��M�����G,A8�?識�%+���Fq��ں��5m8d/��u�D)�$��I�B"~�lu����{�}�+bH�����MD�1.��I�y�DWo?�������d�8w!�S���6-�'M
�UQ]Av�"��Η�cqX�ճ�D)�F8�C���E:=�S�l6ϔ6@�e�)>>Nj���FM:�Y��+������زn�t��S��\���ϝF�RXN�q3��_���7���n�~nZ��E���3'D��C��CA�dɪ�X��<�׹}������=�޾K��`>~�ӟ"��>����A�Wm��0\�.8�PДD�$���XؠZtttx9r)���|ʞI��	)�o�X�t)��������>uL�;s�)\D麞����s���};��������Ľ�vB��g�K�2{Pu_S�|^h��}�n}�U��{���ݿBˬj䒓���6Q[��+�*dy�'�����Q{��Q�x��^r�XE����m�֭��<-Ԅ��zFRP�0�I�jMFԤe⚒��N�&����@Ȟ�_|��0�z19���(��jl������J�����<wXD�ʅq��!���{v=���磡q6Z��A{Gδ�A5��Jd���X�8����C����t�̯�Z����3A����af_9x�<�^9%�ٓWrN�9+�
c�*����<{�O��hYFQҡ�D��a^��XUo`���c��"KBs��Ѓ�Vԡe�2�[�j��%���:�긆��8u�0d�Ĝ�*X�ܲ����C�l!^S�`���:����Ǆ�����fX��S�i�]�|s�)�����6#�#����`:~8zG��4� ꖤ]��"��0���غi5��c�s���C���Dץ	HZ
h�B�$'p�W�S�*�A4O�.�	�Yݲy7^��i2aP4�w��>�g���th�b��W]�\�]ħ>���%�']���2�Ie��4�U�u$+t����&�ZB�<?�/}�۸84��d`�D�� �J���:቙�PKY|�SAf���0�*B��x2D5el�yQ�lrB��J�Y&��O����,�/ӑ2�[�R���?�7�_C.��>�8�{�Xr����J�E�ă�z�Z���}w�	�m�.w	�$��֣�:�W�6��h��'�Jl�b��������%��Sشe3���oal,��z�H�t�V���Gz"�冝�!,L��iJQ��g�{t��[�օ�����3g΀�x�4#7Ţ�`0ȀE8El޼_��W����G���s� �vU��؀�[x:9�����GEޖ0k�<��>|�?C����`�Mp�����@���@�ڂ]Ăٵظ|j�>$���8E�UU �#�q�K˜F����vASQr�������|~�D����s�2�{��|��j����I�j���R
]����0$��`�]��px�WFS���\��>�^,���}~YFe}�p-��_��@��<~�����n!�Y�	]wYߖ˦�̯��&̪o���v�G�v@�TFFR2����l_�'����7��JlYT�����Ku�f��:��K��k7sȯ�
:qB(fr(S,Z8�='����L�>$��[���XZ��5V6���t��a�`��"�����R��Ǣe�L������)Qʎ����O��9�P�e8(�Vs�>d����d����=(8a�F�S��aL$�p%�D:��ʾbg����"�{n��AD��%X�2|�r�R �Q�i#,�5��^��[�v�$�BQ��|o'���@2*
�QJÚě���X�\�]X�<$�ƢY/zF]L�B�l��)N6v���a����n �G �!�2)$�:&{��T[�w�};�~�V��&�����'�,^Y���%�IK"$��4mY\���BtL�{�_e#��tr �`�.Q���r&���_�Z��Ɯ���'G�Q[�`������ ��*���3L��ƶ��L���|��<5���I]H>�7�|M�v��������\�@��bf���̫G���=wކ��
L������W�6}�g"�ͳ����<�';v�xA����	j���S��-[���#����D��t^2�t�� 72r+�@�X(�����8�ݯ3Ph���E�SSS���n��������< ]O��M�̲�*#Q��uk��/����{��Qq���ϧ�z�b���IM&�̝���9���y��3����n�_���ӷa��,��%Zl��LW<�q)�`���s�0��
�Az�����f����k��҅/���/������K�΋���8\Ep�dn��z�%K����'�TX�<���ZQ7g-�{���9K�������P$L��X5?;Ջ;n،��u3&{����N��}1�v$�}�}�_l�� e!	�A����z
�i��"��+�@�D��ǟ��֢B�աc��='�q<c�[�ۊ�ִ��Sذ�?6y~E��L^�
��D/Y�f6�����3����(���|c���{�"x�R�A�����W4aE��5�C�^@z��sJ����1H�j,Y�	��<����5>pZ}.��Q<�����aPv�k�P����R	�MMHf�8y��#y(�F����A���I>(z��m��2
�8w�ǘ�J҅ɴШ��+X��� -\-�-QrT�y
9V�-�05�?zϝ�����c������|�(�~�j��cx��qێkq�f��jψ����g�´\�JgR�K�r���y5<R��)������}p�8
�g+'?L�y�5���y'�$�;o��AJ��^�� �9|�HRwY���$��0�E,�H�E!>����O�4D�����d8P�j�J�hT��o>�Q�9��[!J�f��p"6�@���,�ye��jj�IpO����Y(�YAM;��=G�Fww7�m\�!�d��1:�ۅG�9�_���R(b1�HHCCuA�ě�ۊ%M��4�UPT?G�q��Yvg�;QY���ZTWWcɢ�hn~�A�sb�ÿ��D���⾟ޏd2��:G��	�e +/R��1_6& �9��e�e�i�&��v_��Ç�`Aۥ?y��^j<��:^�"��M���5�W�[�������у���V\�t��S쮾�jؔ�S�!Q�@ee��cxv�A���{��%�����-��9 
�2�.���J��9H�ʢ�*�
CE |V�*��r�z�+�x�[�x~�{{���\.�\1���e�(�)/Hży-��>��v�4<��CHf�pu{��EE�2t�L�B��K�� O������Y4��+���7���p�����EeU=S��l�jl���,z��m/���#="��eMAB�)�U�v��#h��Gm}�,Y���.�������`,�Á�QtM���3 ��)lY��M�_����L^x�=�^'ef��*p���p	e��5B(H>���w������8�#d�p��F�oT��%��`:[���e�*|���lD��Ũn\���k�g����5���,�:�#��ېiY0mz8�XEB600�ƹ�#I�Ⱥ�>���¶hE�Vy�Uס�(����cxL�������^���c�X7W�8R�H64�B%��G�'��-���#�F��C��w/ 
�'r��W>�ۖW��teM��I��?�]����AOx��54ͪ�g?�^̥� $p�c�_A�X0P|
�Q�j#�u�M�uQ�ԝ19m͋��ce��݃��AND���h����▹�����"uL���ç����a$�@�W{��rlH���8p
Y|�}����X�X�.���­7߄�D�q���V�iUx9,�'p20!} ��Y;8��{��=��f��x�B=���������Y��pJ9Ȣ��� jc:�߲�A������黄Gclb��b�ܹL��L`���hl���nwg�8x�0��S���p��	�����r� ��/�^Q�	�I�A�xٙ�B�xU⟭[���u�o�����>�}��ȑ#VH �͛D_�0M ,,ZԂ�~������k���$L���y�V��%�Yee����{��?���"�_    IDATY�����D i,L��M�,r�%d�Z����\3�_�� 8��h W.Òs�0�w�y����鳧X�O����	STM����a(A� l;M�q�b��z!x��8j�{�00��j�a�2kI�~�j��
A�#�m+��{ߎR����
?��1o�z$Z^�����������y���'�&��a�H ?�޷Q�@ݬF�۲9���v�C���)	i'�������?Ǜo�[����㕫_�B���35󉯗
�,M��x3��ګ���`�pJ%(�0��d���ntOQ�N��Y\�r6��(_@_�Y���Yd��b󵷣fދ݇^�ʍ����ba�SH�~�h���s�́�UdKӜ�L�)�>^�H���O�F礅����kA!|~E��Cf����TY8f�]�Ԋ�3�P� 95Ѵ�t#�	��ִR� �)��?�n���륶ɒX�0�'{��}�$F�6�(*���>�ź$�����5O�ÞC�p��YʔD퇬���J"�S��7���bV���	��(�����O�F�j.����Y��лގM-Q��D�09����^\�ť�!�"](a2W`��)��P���V�7^�:���1��(>���ƹ�Q,с,��)d���
�����Nt����5��I$"!|���;�]bjj�*�j���0�pȣI��*Ө�E�"Q��3���g�pCͺIådg.ap� �!���f���5��¦*\�i%�#~4���`�]�o�����0:>�M7��n���&�h�P S����ۏ������#W(��B���r����D��y��s����`�c��ںj�k�˓�'ePC�p��2���(ؓ���r]t������h�U�~��ض�j��ϊ3�[�}D�:w�n��&,]�����rʜ���_<��#!e��M�8l�Q�����t�?���3iJ!ņ�K�:`�����d�Z�w��ޗ��g�`� FƆ
�0����Lh"6>1���q4�7ï�����5t�_�ai*ں��1C��b��z�'X�� dYbS���@s���n܀w��j�9�C��QSW�peZ�m�y}��������{�BX% �|������*�^� �˗���{ ��z�nSv)Q�>�+����VlX�4@^zZ�K��0���
��+0@^�ghf��K+p�B����:�#�d	@~��At��PT|l���L�Z[��������%�&�fR��Z�;��n��K^��,;zJ�ؚ(7?��7!,Jr'W��k��H.����Y*\��(Ύ�8�=�q[A�R�)��.Cu�����/!��h�*�$�,���v�Z0������r8��)��Qܸm>��wB���������O��>��A�[X�O��;aP���h	kRˍo%�_Q� d�K��D����R6���o�-x��a'����?~?{�i����r|���͛� �L�ϫ�J��t�H�P�UH�0B$�%���XE��WÆ���0�b~|���˖�_~�#����P�0e\��dA�LG��g�	w߾�.�Ţ���[W	Cq�v�Jh���sgP]W��[p���|��8M�\��Et�~�hV]=S�H�:84���Q>r��J�PFA�18Y��D�ȔX��K��8IvUUa	ɂ[��6��C�h�M�H�Q[U���Ztu��\*���(y5�U�Y"kg�@	��b�ls½�Y�z�B"tJ�7y;4頩��ŋYkC�WS�clWK�+�V����@��u�w0�:p� ��v_�.�u(2e����]U����J����P�x.W e�,\����t�x�E��b	S��'RH�� \�W����&�<UF@ �;��6%2L(n	�b���ݺ	~��e˖�7�Y�p��e�|&lͽj��o�����71ə7��
6�z(6L��ٶ��ۍ��n��ʘ��y.�>ER�P� ʶ�P8�r��7��]1���w`����8,��xe=��9��~^ϯ���i���%���]H�P$�}�D�!�#!,]�'N��D��@�i;�4*�'�!Utp��n��Ջ��z՚����4s���
��H������k�'�Z�H86±�2�t⡽�1�u� q��+����J� �;?΍Y�RʱN�w}�e��
�6A[!��g�&F qB��/��E#np��XD��g�I�kGZ1�g��)E��A33�����\;�����w����уө�:˳��O����w,��I��[��~�/�..I�E!�;݃�~���ZBA�6F�� $br�l]��w�>
j���%����Kg��OQ��P�8�I̝[�m[�#
"g���A����~��G���ve (@׿��<I��\�V�C�����od�'�?���7��r$�@&��g�,Y� �=�$ �9Y"`T�ae���ֆ�]�Tƶ��P�DEP��%��m�ͼ]�p�Tuu�O��"��D��]U���<�CA������K/��l�ij��ى��<ʖ��d?�'�(9�BS���GF
��	4VGRJ���� ��W�`o���G�i�
]�|I�R��%����2(�����q���y-(�����s�V�,li�A)�TSP1�V�p��e�������X�N�� ���2 �G.���T.M#��P����I�8_#��� J�́�rHT,����(X�h>[גEv2Y�#iMe084����H�,�9�Hԫ%��S���Î�Dv!���0k���������
K�,�򕫽@K��q]�+"l�K�E@,��bdhػ7)$G�@�А+���ۍSmm�8Џɂ�Ф��D	�b 4��΀��Id�k�����ބ{޸ǟz�}]�����������?�^����K��2�k§�:��ߏ��~466 \�Ơ�됵C(������M��o��7���5k�����p�g��Y����yZfv꿫�Ϝ�*L ���SE����đ$mҮ�uQ�\��K�e,���{s
�,P*��
Djp�=�{����y��6$;��Ӈ�s�<O˄f�8�"@�TB.[�#��(D|!9���'.!%|(:��0���Q곕Ů�}��t~8)�@n@Ǧ��'T[6P"Ṭ�uT�v�ly���E����k�Ԅ��š�C��g�kNtU�u��O} �tI�6�(�����v�c�27[���3!7$I���@Τ�����!f���%ǅA���x����F�����\,��-��p��6(�VR/��@0I��S]�V���[.����02<X
�Pv1�t�h���-aɂF�r��`�%�MD������C��WS��+O��e�D�I��Ȥ��lٴ���ٳg#��G�O~v?dE�d�~�N��u�E���@�JP}D�PWE@*�"��85��#�2n^S)����~�D*9�ʊ(�G	~}===�:W��4����j�%��9|P���}x�2OEH����͘��D����)9��d�0�)Zu�D��^{-��ĉ,�'@C�/�?LM{1&kj���[7t̞یB�5$J���e�R����o`fIy�a���m(�eh�0_ӎp�f�� do�Q�l��h�@Rh�G�_E�ٓX0�-s�ફ��5���5�� �_��YU[���N�>D�sp(x��=�T�D<˵p�������Չ����)�!���� ��#����D<�CD�ė>�v,����ܓl3�BX��
���?����ٿ��f�:E!7	U�a�2�\
'��b'�܏���~uMMh�ꇣG0i��Y��݃I�p���q��'Gq��
�oS����T�7+0�P��f*��w����hr�Rt?&r���R�M��5öQ�:ض�+�\,�ӡ�����|&��;�[�a�?���c��!�t�̜�c��q�,� �o55�,;-Q���h(	?��<r*�G�t�
�aJ27Y�)��(N�c�Ͼ�u���60&$�Fe���z�9[b��9��\�$�*S%��Q\�q9>���cUT�.��x�X���08U䜏[�Z�?��nN�̍K�e��=��?������
���$\6-�%R�r2h`A�$��E�aAt� D)�����*=�z�hR̩��근Ae ��	v����j�e��]� t"Q6������6e/�LɡF��mAi$�a���&�A	�σ(N�&�GCM���/K�G�Vq>��Q�M�����񤧷��:U��34d�R|N��(�����G��dq�R?��)����� �� m\t����	̟]�Y\8w��:TW�.aF"ynU^�=)6�VF5� �.�P�S0Y풛���G��
&�u�a���9|P���N�H7Q,X�@��'�|>LP���Ei�`H� ׃�w��z+����t4>�M�
�`��.J�)������̚Ո��Db1��&�4���ĵ�H$PYU�K=c�W�"gZ8s�%���'tj�3�C�J��)A�Ҙ]�o������چ�ߏ������xN�<��D5f�S��l���	��v±�bG�0V�]b���}���8z�F�%��̹Z��_�Di�?- 	-t?��ÝhCf��]₉Y�|�m��^��Ы�d��Qahҩqh:��
���#�����������ݏ��,U�(��8�6����a������7AsKغ|Ɔ��r�g��W����+����c������C���
�9֎�g.1 )HԒQ��.X���4a%�1��	Iv8����������r�RC�"�!�,&G{p��^^�We��h$X��u��Ua�AX�9x�L
;_��@Yѹq����Z������X_�Jm}CbqS=Kl�[b�T?[�*��C)��NͿ
�[��Ǜ�ۄ������-����g�����A��ۮ\������8�#��������
X$�v�!&}��Y��dA���R~���%�B0ǥ$
�B&Ji��X� �����c�W��.��ԕr�LYDi��ە��z�s/�[x*.�9�G�ƜhO9(r	A���m�R	��Ϡ�"�������ɩi��`k�x$�zʇHe<pb�������7��h���g�ۏ�%�p��<F�9�MP�5؂D�*Me@A�F�DE����*G�z8�¤�L�\4���%����h�$@ A�eXf��6]�������`�A`��S�=G�g�m�Ώp���Y��w�},(�e2�G���<Š�M'h�@� �N����x�@W�h
C
��%�����8���?�	��(&�)�
M2h��"M;z�_�j���Lg����Q*Z��4e���D�p0�����&�`�'�zY>��'?�G�r�Z���6o��0�l�A�}�ͳYl?16�������3�\�T�,�'!|Z/vch����2��%�dB�A�A�&[HDU��8��ʇ1Ҷ��^�cU�,�~����9�r>�^�mO���rʳ㥴'QFP�qx�^��1U�7�|�EU�5�������}��܂7\w�}���<73�z}U`���:�3G���َ6Q�˼�M���б���;�v�EYg��Q����s�f��s���a|� l�d��C�ܥ�z��!/���d�a�����x/���a���M+����iBd�}�����(g��#x����	ٽ�����[�#��65�R�Ȕh��K��+��N���c�U���A�JW���Z6!���7���V���1���=g���_�)+�T̎_����A�i�I��w}���Ov�EHD})��Ze�pM�M�Kc�/(�D�X��.�4�3����]��S�|H��0�� !�{��� 7���Z�'2���
85���I��	�H�@�~�-Te���'?�>�U���a4VU���A͇��An��%q2�����zbn��8<� �@�B� �MMș6?��W^�ǞڅξAN~O�@���8�΁��F�8�� �J���?�,
ԣ������4��\{��*QZ����	۩�N������JTh�A�wj{;��s��7\���_�"b�g3,��NH,N9 P�͛Ǵ��;w2�#�M$hr����u$��e� A)�ZNL%Q�4C�d+LxQF![���*��4F��&l\��W�hڜ�!�	Ӆ�.O?���G炂:IW��(��Q[Ľ�v�}��u�M8��L���7����R�C~,h��`8�'�z���l_5�����N��l��L Z3{��@�D��#S&�`�)璄�A�������p������ѧa��MԠ~�*��t����o<�sc�bj�Ѱ�\)�Sˠ� ?5�]�<�Y<ۮ؊��Iց��2�@=�"��e �cv�,�T	[W��#3_�3x-W`���Z>�3��[W� �-	H���#�)K��z	;��Ř)�D_���/fq͊&�oR�q^�y Bڋ�Y`���q���a��o�S��_����ρ���w�Μ<��U*���#�s�I/,�S�����)�<�)^�4��A�fY73x���+��?'��Bl��n�x#J��+�Z,l�W�-��?A����ڸ��Ľ�` ��O�/~�Ș2;Z͎J�Ɨ�����6��	���?ƔK $��h�&ʩ`[ޘ�r�*^"6����m&Y���dN }�=������#�t\pd�]j�mɛ:���2Պ)Z2Qr�f�p��9�ܑ�N	��Ļ�!��������dN3�����!�>�οC���>��0��O+�&H���Aִ؞x��xr�^�eK|Ț�M�tcԬ;H�	�W1� �@��R%�ã^	����Ѱ����ҊCVt�ehT��Y&TUF"�U�db�y�b
m�&C� ���hU�_=;\}�;�A]uOvHkE��ʕ���EO"sr�":	�	�E�(X����(X4����|�t���������ih���SV�5!tr]Gٶ��TPҽi�yW�3�kI�O1-2h��A��1Ō�B�U*��_�iH�櫷���	l[��m�LY��k��ю�����44����Μk���%��0��U&��
�Ϗ��14,X��'N�|�
n�y��ue? 霻BTQ2>��m��m�/�w��d�HT7�q�&T/ya��K��y5no�}��e��<EU�'�-�z�18����#W,�� ɼ=�Y�@8�U�5HF[׾<�N�ƚ���L~�
� �߶b3�MW�L{�(�J�#`
	SE����G�0Q�`�[��]�]�Vϒ��9k��}��k�U�R1���f\w�{!// �j�b"�sqd�S�pA�x�F���r�k�dEICA��f<ur;�k���G�-ׁ�j�>H�I���7��F�.�e��(�6�t7kDY5P�&M�!�*��m��5Q���� �ٴ��Ľ� �t~��|����,��C"����@XFHB2����@���vlrn*�e0P�OM���{����bx�80:,(VSG~��g�o��8�5��A�"m�1������N	��׉�C�l:����i��\�hş���PDk��F�' �IDh�s��p���sP%�x���\p(*��Ӌ�:(a]��'��N_�A0Q�'�;̙d�;�.�r5�2%�{��6�8��!�ɍ,���1�IE��t������Q���Cq)�͂B�N�	�`�Wr{K�+�������<L��,)@u����}>?�~�iTTT��#��=�e+�N400��=�z�IQߦ֩铡q���$�$C(D��1�La͆M�4�흐aD�UH��|����&X�!q i����t7��%���c���T�ៗ�N�p$���|���D�V-B~x �J�$b!?��s�h�o@mu%����c�x�d�L��$�O��J<5��2��h^�?����x��o$������@��b�'#��yq��L���&+��mF���H̽r�{��}kM�����Ѵ��	���8q�����j�j���� ͨ���QU3�p%�a�%nݸa�!A�V    IDAT���`��^�
��</gug����@�"S��:����
�
�N]�XI�	�c�Q)ٸby=�U�X��4Տ���K�F1�E�����O i/�P1;�!�B!	O<�c���#
0 !169�f�'�`/IJZnx�kMa��V Z�"H`O�k	�@j1�g��:VUH҅�)j҂Al��N��F�[�&��+�~���"#9ҋ��Y����p.ʶ�o�x'��^b(�ؼ���Ļ@�ڴH=�t�?��'()ؒ�T2��T�hO�ʜ~v��)�'z�$����	�*8{C�SH1 ��-��.&a�!�$&M?�@.O8Ƃ�M�Ƚ�.k>$jLi5|:\�>�vLH���!0�:���1����]�܂r>���^�D&�4���LSSCM����eҘ�J �Pɂ���p}!<��Dk�.L�-�P��N�ppc���8S�Tg�d��^oBz��xG��i�x]�H�b�<�P�Ś�(a�<tEFU��\q��D��u%�"M�<�_װh�"^����"�n����M0� =��ҵ¹��t��W��<t<��5?%ۂ��#ZY���F,_�P4������݇@0�\��*dUe퉦)�����H��R�'E��8�H
�\F0�Q�Ȧ��g�=��:˳���3}f{�j�ժ�j�E�۸�1%�p�%��$�OK ��)1���WY��{Y��j��v�w=ϙ�q���8`93ץk��3g�y�;�<��܅ȃB:#�8y��(��!��`!"8�lm�8w�F����LM�#��� IBu��!�ɮa�o`@��4A�[=����X�gv�ƶ�G�.˘���0�ϕJ��L���i���-���/����a6	h��-s�"ܺ�z��7w���~/�9�PX�!�\DX���sG�Bss#�[��wf��	=L�Xu��턪�9C���9k�W�����Ww��2�/��LT��1@���}$=����������ι@��S�8Y;��YXҪCHsD�%�˛�<�Po���!���~��'<I2�2��{����� ���Z�n����&'P��ڀ����=��(!]b���S��j���}�Ƣ� �$MGW<&��^�)�ր�"�Pm�"tY� [/���e#>�QJ�0�L�k߽�?��-ݜ����_��'�ъ"Hć���(	QdH�����9�SQ~�wT)6�Er҄H*gqP"Y���`�{�|�}����� ��7L�"-DE���麚���z��\�1U�D�*��cb��Y�������t`��b2p���p�9��<J8��Z���B��y�̠����[ 1�G�eԆ��׃���&�0� z��׷�t�&�0I�`��A��˦}s�V��X2�H�����;[��n���~M�λp(����-yIנ*
;xe2i�[��!�At����TX�]n(`^Z�_�b������4����!W$PA�a@g���?W�HB��f�e�X=DCs����!���E��}���Gk @&7�R	�B_ؤA!k*��H�D��x���;�j�BDC�!�� �<�� �)aN{=�v	^>��AW�\q٥�K�y�?r�e� &����1u�H�ϡ��EW��m�X�z���s{a,� ]��clM�+�lt!jC2bz�h�e+�P�<�P0�9�נe�z��jVſ��d�0 	Gt�#
!�J���}ܝl��@��0&2�k�Q[�U���0�,A��5U �qWw��������N���`�
"t9m�(�ض�xjO/���d��
�pE��X��75���S�l�ą-���.�͜A����F�zA�a<t�`R�Idk��T
��`	�����(Fs2N �%}S"�OA�4p���O+ܒ�Gi����MNy�jj��E�ZO���G:�da8����'kT�����R��|��2�V8>���ֆ�[�z���7����D�bAn��a}ȩ��V���"H�xj��i	 (\�,Z��i��yAX����>�6B�LQ�ؽ�'�
B�ȤG���za�5��&��1����v��hN�>eZ�&�?T�6�I�]Ř�C�D�C�`{��!���W�)�d��X�����C
.ٰ����OpW���!�l�j9~u��'a7ќh$Y����Z.��A��ᡧ�����G�����.�A�3�����JH4�'�(&�� gvXL*;Tӹ�9��QfG0�:+��lF�YT�H���! �6�� �z�:�
?��)�Ƴ�+r7��@x��:[X�^����l�8T�N�&� ������x��z�:�Z���cޢ���$>w��16�"+���|w0�U��]"(����ٴ�"i�h�yCz��	�t��3T�$Y�y��0�{�� ��T��o��t
�l��t��!�<��$���h�$�;A4�(/%�/"S�F�x��I$b�c�2wb�`e�c�D!zA�B]�Ƶ[cI��4�p�s���څWT���V�8�K)�nާ:<�B,��>�:���&�$�0�."^ׁ��9���R �\Ų��Ω��늡z����~y�3�W}�n�>�Q�6񿡄`JQ<��~<��sSv���`%�����/!3�rj�AnM����X��\�_�B쿦�;�E���T��8���?���$D\~�;�PEW���Ǒ�5�D��8N�)�w,O	2HЃ\�+������}sÂ@ ���:�圷z)C���9�0�+#�E�`�
qmDC~���B|�?�ٵ�pb*�u׆�O��s������JX�����Oa�.��#'م+�����tZ��m�P5�Zl�j۾�,���h,�̨SAI�
��K*v=�#,
©ɜ7�.�׻5W}�;9�C	���bP
5i�}&U䐴0�/��t�r�ݯtEG!G!~�_$�
�ܨ�\7�p�*!�	���h�����,��0Av�%ޗG}�����Lb���/�wE�h�8��b۾cPM�@A%�W��ALO�f����
�k�ȦR�T�]�h�W���eS0M%���*`�B�� ��|&ˢi��%Y������X`J"�~A�+�G{���Vu</)��^�������E�����������h��<d
��_"���:ΙۅUk֡��Z �����a���^z�`���cC ��i�=��.H�b��� @N7�I�g�?F�Q���U7\�<�˟bFmKf�DM0��^v	���Y�� �P�&�QI�*`�:-�� -[��,y�I�O����@
5�`	e��u�	��ba��b��`15���Զb��5��i��� H�W*�`�Y((�4:��~�3������Ś����.�4t@�Ȃ�R��Qv���y�� ��Í@�����'�#���/G�ڂ
W�P�x|�Ql�yC9A� ����s�aA����"��(�F 8l�B8�i�hk���K����B����Ϗ��B!dK���c��(X�̒�'�X��`
*~f;L5�����X�=��C���d=�v��k��ObǓaM�U��F���M�m>��v�}8t�uM�(Z��-�ЅR���|��x�ƹ�\c�����ϯ��
ձe�����/3e�&�s��6_|5�Hf��<����Y�K�MD5�e�ICa�(��;z0��i#H��:u�nw��Ul�������{i[���΄D�f9�5a%����ba�?o��Cfr�; �X�t�E�jH���y��Ҳ-D�:>�ɏa��!<x��0�N�_��:$t�G�� ]���(s��,���$�W����#R7�&i:҆��cYl?z;� �<%ҍ�{m�`�$�<*��2:;��y��lGPUp�TkE��7�QΎs�D�4tu�A8c����~� 93��;8��4�f�~�8dYK�,;1r�b7).-^���N@W5����8�^Q�m�������A���&r�<�٩�A�,/��EK�p�R>�H�3g�ǟ��	���.v�"M>�7�<�M���=4���O���䀁�'ZX��:V)X&���|���`FC�\���3pٖ���g�D8L�U6�r��늬�:�,[ �9��ptݠ�Q�p�.	85��Oي�����)(�H&&�"a!���&�mY�Fi
�]@}S��F|��{����N{�b
���&���JC	�>� fw�C���Z�o��hC�+�VсcX���������.�1G���yc���^��F��ɣ^*�eq���(
!<��{����Dtl4(6/i���U�Ǐ#?��T!�*�&���[*�f̞��y�m?�u��y�#�FN��у`��p�2\�\�B�����Z�w��W@�	IS�)�a��1􏑽��� ��"j��-�s�A\�~)�ά�X�7+���6�;���}hl��q�5N� ��������U��='Μ!.�%�×��T���%���/�q94f{K�^�D�Bd�~"9i!�h4M����㦦���a�0��Ȩon���+`�$�6���gn���z&�l���3��[�㩍���4r��K)� a��~��ًhG��0P�g`��L%���(��1�ݟ�Ԁ�*!��	<��/��C�b~[����Q,ݷ�;����rV��n���>�W�]��Pde���(z"�L`���91c@ (��О�3�׀��X�5�]���n@"@��c4�f�)?��E��Pk�Y�Ʀf�����c���`�T:������Q������V��DB�s�4�~&�"I�cR�4�e˖��6��[�2P������y���N���`Y�~=z�N�kV�T�.�̓@�lr��X�p�/\�%�W��k��������v쁬Qދ��;Q�xl�NG�V� ���o&i����N�+
����K/ڄ_�w�l�[֯Œ�ntw�Ğ];P[�Q�sv5�ϧ������(�G�Iҧ�]`*����$��i ��%�aS~��^O�y�����Үn|�:�#�U���s1o�:�7��ל?ҥ�u��|�WH�r�c������V��D��Ȗ,�%�Ա 5�3٣�,��y
'�i����}��Lu��]F�����r����5Gz�y�\Nن%1�'wţ;Nbʦ�iL��[:�j],������@�B�: �TUG(V�Y�`Ɯ��V�n�9/w҃n`��!�yy�_,�%�k0�
 ��t����f4v��?zV�)+ Gm��c� 
���բT7Ȓ]�0�)��7����y5����T֛� cY����}��%��01:�rn
�lـ���~M��GNC�[[���Ɲ����E���LoZ�����׌�ضҋ�̃�A�P�P��C1���,P2I)��`8'��zg=\U��*�Q�{�� r���,�2�L���[n��X#�hʔ�bP�o�Jz/�P�e#@ŧi��.M���r�M0Z�����!�
�%��E]}>�?ů�9^|�A,�j�goyw@z���Z�,�Q#�A'�
|%Џu����8��L���=C8P ����p\Z[�C��瞅��:�7��^����G�r�o�����oy���n݊U����C>�g��P�N��O���_x�y��#M��GA d�
�������hX�p����ִ~������r��F$���~#N�<�ݻ�2(!���o��er ���8��W u@Đ~e���ꚃ��CV�H�7b2�ÿ�}^�}�m�mj5Q�O:�� �
 _Kê\)��D��@H�S�����,�����ƍ���[1����*�EBhi�����(��4H ���7C � �$�I�e̠sDCy��c;^��G�� �1����h��w�4�Df5x���P�Ͷ�3�,Â��7�~ݮ7�Wг�E��q ��!��P�e��{�J� �@�B�s�j[碦��"A��&�� ٸ�
@΢S^��7�T/No�Rݝ?�P!u@<�eA����؋��mG�v(��UD�)���X֪c��Tc���ȮA�,r��Y6B2Qz�ͭXs���|z��>�yN/����Da8d)jXP]�����32�B��.�̞����)�^y7S����@�5���]�CH� �"��Rj����C��1���;6��j�Oy���oEm].�p3�?w=.��)aa��5�˕���)\s�{a�:��f���H"��`~�U��7:��lj>�/y<���$��2��� }�k��L��>�O�op��˅c����q��;~��^��SQW��w]��\�V891�I��Y�������� Җ�`�E09BG�"�%n1�h@B�5�ͯ�o�5�8��4>��/`tdҟ@b'"*,=��p,�|6���>�g���߆��aQG�w���8s���H�᰻���|I�B��!��H�Cx��`8%��ϼ��G�P�#(�*�����B$��Y(��bM��f 71M0pϝw`��ů�ޟ:u��������[�p�>v��r����ߺ7�~y������k�5�\�[n����u�X�zH��m�t���sr�:q���4�����Z�
Ǐ�ľ}�xΒ=/��)5���;w����$w`H�Bb{�аvDEM}-���J�75�#J��cl"�ށa����P4l2�b�/���p��Ҿ������/DUc����@�9́����Cd#�k.>q���� .�r$-v�b�P���4?ѝ�%��
����Ɇ���ĎC�1aX��&(zD�<�\JC�L� s�\u�h�>�U̚��Wl��P��]w���)�X����n� ;]7I�MM���qD(�(��oF R5����J\KĚUU
���]���y� �l>{�}�G�H�	o*��5 ����m�����1e�():L#��]�Ⱥ�VtƠ[�8��s,P�4H�Ä����$[ۚ������1��&��	12=����3�Bjr{vo�cDXL��JZu&���J�J��{�m�������J-��h�$��$�4�MJ0�S��b�N@X�<��(n��r�Ňߋ%-	�����x"w�	�l��cӲ�1��(�G�e�����m?�}韾���Id�6\QC��v)���	<��/�r:96捧���?߉��
)�+Ȉ���d)��R�M4D�؟ 7\{5��a�xɋ�����k������`>�����w��.Y�3��Nغ��������F���=H:AF,�@rj�ذz1��r.6���H�����_���A�$X8m6�B2�
�<�Ē���؇އ���?��� ���<��E��c�;�6��c;��ӸX�@bt?O���A)���p�����9OC��+Z0�K��F�}
.$W'kV.��P+�o��q���u��=uһ�߂"*���Ngq�E[p�[^so8��������8�;�||�ӟ��@z�1 �3Y(��w�"]�951lذ��)�y�!�pBz�֭O��i�kb�V�^���	��O&y{�I��\O��}����F|�3�4��	��5س�0F&�x��at|�<�|p�9�O������D!~G�U�j*<��0�e���.�&C�m%5������EW[���Rd�I��P7�rPx\h?�̀�gUP�$9�1�K�tw�N�`� �Je�]#)��'�0,�AQ&
�*�� MQ����Y�!��X�t��!���u�X��L��0 Q�d�f� I�TU��F&9Ǝdy���hB��������H咋�K_Z�Y<��]����5U �{W��o�8��� �*RU�i@�~�9e5 ��C�-�%3�z�����Q?��UFX� Z.g&Dd�b0�� H�������D�Z����z�i�ɥ �%�i�����0��)NZE����B�(>�-b*_@׼�5���?�qC��գ$���@'N�0 1Li@X��s�CA�� ?5�����^X    IDAT�
_���^�n�f�YM>%k��`�[:�Q8V��CGO�����>���Hg��C���B�-5��o���0���qx��[��!���=ޓ�lC�h�*{k��P�q������9��]��Τ=K� ���ԭ���/�+��e̛Y����w���M��3Iv��Z+��;��:|Omۅ��z8I�T�a�-����?�u��%�@4���d����c����E�(ħq=�,2����,�����]x���p|�6�D5���-h�K`�� �r�x8��2|T�JӰ��x�*sW���R ��'�����0�(�
�($9����1=@չ8�d�8��eă"���ױ���5������ߺ�;,�H��
�F��݌+���5����zO�Ʈ]����x�R����d� ��(�4> ��ۧs�f�457��.��H$�E��ӧ�}�N�B�E�+W.G]]=� �X(���tl۫2MK�(���nz'6�w>FǓl}��	�M�𫭿�ɓ���nW���X��~�f�2},����!�A?Nx/���0���nN�+�����7\}-S)���!��'2 a�� A��|Q�d��Ͼ��8ufä�1�g= J ˦y�1���-5*�"6-mÜQ��[�	K7l���9������+�V)��������2"����]VA1�L!Y4�)Xb �e�T<^�r�ƪeՔ��.s�z���T��?��-��#p���KrL�� B!�g��į��@�dEYE��E�h����Xծ`���� �{���D��lhU���B�dB:�����kBB�6���`�E�A�3C<��s�2'��.�THcrt���F��1��pH��c5��kz���Hf�蜷��6|�'��hId R���ӟŉ�A(� gQP�YÂĹ�S�H��)�N���%�{�]��P<�=��)?<0��8F29�觏��_��x�T�h��J.0�"4�E n��w��?x���\֣��Г����k����:5��ʎ���1�+n�>��o"R?y[d�)+7������r,��sb"�u����/�)y(�a'r���'8��/ݚ �(y�ؾ��N���{_���8�3�z� ���N�r�k�1X6����-���;�o�Ө�x�;�EKM��'X�P:�'�V�S{��c����]�*Щ��I ��ޑI<�s?���0Ţ�|Ʌ��p$�s0������ǡ]/a��F<�п�ֵ����{_��Y���؂xmҙn��F�]��5�?|�G� �BK�/ç>�)�楬�O!�a�\hO�B*��\d��46գ�������'���C�P*,H�N��K8���CL�"g2&�B��7$B�בf�(Xo�;�z�9Hg�(Y�<�3����~�9p��X�a���!_��]Ô1_{3�� D���$p�Ѐ�y%v�]��x%l\�A�;7���bQ��ƛ048�,1��*��(�K�G�~LU4��VTZ@���;8�������d��dN�� �p�2����\ԅ���å�b�V>�YVc�9[ ׽�vw_�_�]�L��J�)���d�|���h8�ft�s�+�1U0Pv5�J�B����p��✵����;Y�Xu��#P o�\=��o�:�M����
����w
��q=�y2%�,޲rV��XԪA��q��a8�� �)�P<QZդ��N@�m0!���c	�5�pr1�K��A+�d-K4rU���b�C}���R�хC�{*��]�_�Rw��NwE�E�r1c�<�uM����`�(0�V�p�/�����Ũ ��!�^M���g�:��g�����5��g�	:��Iz����.,�NzK[k�[�y��ݻ�R� "%�I��������X��������U3�)񤷢�׏��=��MԢ3"��=����V�RR��Ó~Ai�Q�q�%��O�� �! ;�fKZ�%����^@��L�v�8��> �L<�dbAsB��_���g��g�ę�4\Y�.�]�,���	�����g�o?s�����3�BmX�;�v9:ۛ�{�2�$�j��ȗM��SOb}�r1X��k?� &�WZ��2Y0���I�D��p ٳ�eL(ܵXS b^W'�#��h��W��wX��[8�;�͞5����~���W��h��ި�o��̍7݄�+^�سw�GnU�>�(
e6nb "��tH���Nw�t@h��C�;F����6	���,R�D�P��[,���̙â���	��A��v`�-�Ԑ���ukp�uף��S)J5��g�a8|G��b��(�!sv�r���ȟf`ɘ�����e�ٜ50�[�K5�(������S�| F&�\��_����D�S�i��|��L�B�ˆ��p�OAgPd�l�B 0@Ͽg��Yᡧ��h�����l+E�+Yp�h,D4Q�p��.��"�Ag�2,���M+���ѿ�={3���=�S��=�ٶ�ϥ�������!�|O'Q���)C���A�Xw�s�nMU�f��c�Ì@����꧜%#�s�>��\ۃa��N���0�s`RR�]f r��N�Z>3������Ü�&�iA�=�D��<�� d���P{B�Pv��e��8e��8Z�!)��*����q���	\��B�G@ �|t�pV�/�����a<��H��߹��ȸ,�	3��Q�S�J�ɹ�m!FK�L��P�\29�9u5!���_���/ۂ�+�sj7Q�N��ᑧ���<�h��R������#Ԙ�b�4ED1��Q�@�
�5���u���ߍ9�u��7U�f%��N���+����N����S<��~�C�DQ.�	 `d��P�&[x�5��#��t��H_��ҩ,���4�6��ˎשK¿l��}�� ^ۂ��C8��1H"T���.���N9�y����W�;�y�_x
�g`����5���z8]\S$$�Y�-ink�"����m��0����d�����)_g���5�G?{y���H�M��9G ���Cs��j�D��Mk�bV[36�Y�I�M��#����B����Ba�^\v�k�z{{<r������pɥW����`J�IT�8~�x��@�g�X�o�e��A�����,��?66��7�#!�,*��g�LPW��T� �#�]k׮�o��r�µ�����n�ds<� �ӢUm����\��5>H�X�T^ ���ȎX6dI�C�ϔzo�lJ��_���s���%PH%y����`h��-��Q� ����4X��(<&�|�QD,�`|2!³;vr �+Őʹ��qX�����`�4Ն�X>3�����H�4���y�\�pՆ�w�yr�^���k�9�4sPd��t�?�s,^��-�'�Y������3 �I�y��?�J�:Kn���|�@��OJu��x#���Q�hZ�lD{���O�����H(J*������d&6+fG�'1Գv��h@�DV����	�
L �:���+���CE;!��Q�OŨa���r,^Ae �K*<�$�D'� pNk����0�sdZ�P,ۘJgѽh�X-~���HZ

H m��3bbx$�y�>önnF�ܹOe@�Q,��ʒ�1�-�s���)����p�w���H�X#!�d�,.iE^F@�LQnMC1�GkKFG`�3�>��?�5���N���y	��_}�ZMf���x����N"�܎"uB:
���T�� �BN)� J��7��ų@y�ż�E�H��Գ4A؛������&�Ҹ�_��j�z�޽9�Sb�+@ N�aCVdȲ����Y-\��ؿ�wo�$���(fu�c��4<�ٝ3�=o>g�D��y�UѶWE��=��/����>����3#���9�/�]<��TE[D�\�a�5��Jh����"
jB
���"^�]6T��Ƒͥ�ӇD6�c0@A���AZ�K/}�k�������}�W�r�t�*���I�̧s@�w
*nX��Ɔ:"�N��/�\IJ��Z>�ɟ�,(���O=�k/x��.[����J$��)X����&l�|>f�쀨Xce�">��O���0d=����\� �Ojw}�!w@D�n���`����kE�F�ܹJI4G�l�(��9���~�\��d'�9�q��(���F�,��G�hmi��G8ES�J�e�쫋E���b�{�#�oj�Ï?�S����*C�l��:��(;r5�t��n����c��^D"u�r���κ�z������!����4���D�ģ=�U+V���Lf��� �Re3�ښ45&خ{ݺ�����ݮ��|��@��s����#p���˖h5҄�(�:^:܇{߅ђ�� ���n��bYG ��4��q���K DW!�.�d�6�
m=����.?uHd�]�Ӣ��BEe.�"[��pPGH�T*3�E��Z��dB�R��r"W{����q�]�j�?yx+R�����ĉ���������!\_���V����
V��A�N`v�2�ø��װ ��g����"��'��D@�q�g'n�ը@�D1R`�6� J�4D�Cg[=�cg�g１ݷ��k�T��!�,�|�ݺ���:�݇N ]�!jZ�Rr�:G�N`Ig���hB(����ى��Ly�NRwwwE- ��b����Q0l���p޹���3O�H��u����o�t8HN���EwG���������s
۱Z��ف��>���`��y�9{�ε�[���ޣ��P�2S��=�u���Hϱ�^1�����x�ɧ����p�=�d�jc�)����p>�\�mA�Ɔ�lI7���o�`�q,�ׅMMHD�ŷ�s;2��̟?�O+_���U 2��;x� ��w�ib�hw|�{h���-�+�s���t�G����ڵ��.4Gi�Ӄ� ė-[���.�����022�s6�4��>U�4�TDݑ��ź� (:[[����N���s�l�������K��I�x^тT ���<�D��ȶԒ���"<���F�=�'�?#\w�5�9��!��0
y,_��;J��*2�^s�=3pԓUu�4Ms�������~t��&��s�2EґbK�Y��*9�V���R_BL11�Y�{޶#�� ��" 3��){}��g��R#�<Q��0���F^h��#�g�܃5��� � ���D�5u�B�H}]�a(��M��a��Gu�#���@�����Y�o�898�M���9ĭa�a�:1���؍3yY{�v�:k�bv]u��(�#=-Y`��)T�h-J@�D�I�ȩȔA4/���\؆������.fD���f���]r[��J~z3=<��=IC�$M��}�����ʵ�@	'p�?G�$k1RTП14Y�*�l�J�:*Z<%�qb�KT0��H�B�GcF(;�v����4$��Jh�Pr ):l���
u#pD\Zav���p8�y����IHaS(�� ����&C����2<W�4�Rف!�� <Q�|
��{"��QR1�5V�~�@Wi�yh� װ8L��uc���q�oT�N��ɢ8�����ph�L0 ��O� 1��6��]�50���^�O������#�+�GI��*cŲ嘹h�05��H3A����nP�(i�$��>%�V��t��1==��'�~b0�{��?���z��,C��Q(�0J%�#a�$�V�Q�3�P�  � �J����X�A��͛7c�ʕ�=���C��i�<�y���~ $�L%|%ɝ�;;F� ��1ѕt,X� s�gcjb�����$�;�t3g�<ԩ��F��Ԅ#G�`��"	p��r0�ЙN% �6m���6CV�=������N��r�mCs��P$w�\���k�b%�n��ţM�~!��
~8�MᢒU�ŊU���O~?��_��Rˋt�7��_��&GNy5ͳ�S�^�H�N�G�!r<�����:�����E��w��L���K/����P�z�Hr �EI�Q�D����X���=�T	+VoĬ� ���Co�K~jt�G��F�D}"���^4���N���_>����1�+��U�m�Cٍ���a,Y��Ẇed�q��j�f������@������#p�o�i�E���~��i���]�]K;�~I�B�8�3�]��Dt)�TP��nI
P
J�4烄�N�t���+�6�皜@�Q.[`��i��O�vY ͎C$Nh���~vm�b�k�|s�χ+��ճۑ,	({1d� �pf� I$��p6Uyj"���K�q�FBr�?N�w�Q5������l�S�U-�S��������-��P��3��������+"D���}E��l�>u�cH�bĨ���*)׼�a�c�,갈�!*M��1���!ςB�"�E^��0=��ThE��p@G1�Ī��pl�>�GF �,%>������P%��93��C?��F]���~ͣ��&he��e����c�J'�F�[�9z{{����i�ӣA��qJd&����0��⥗��'~���"c8�B���9DE�.�(�& ��H@D[s�k�HN��*���G��fX�N4'���k1�?�Z��5��===w+�H��z QQy_}�Z�v���Y�l aݺu�ꚅ�^܆���<�:��&�c?���6y��ކ��><�䓰���C�0w
��}�%�bŚ�gvua<��{���C)y�'+N$��E� O�)De�]�E���N��dA�"z(�P3[�~�2���"V�X���0 ���>�ʽu���G��4�u��e0�ϡ1 �*+Pe	�����?{�����܁g^؅�΅��@��`���h���B�p� 0#n��ބ��>�,b��e���<Z����y�)${=�H�#!�w�"��T�ݏ�������"��7�#�(Ɠ���҅�pκ���Ъ5��pc���r�_�7�i���k�9��K%.�(�� ��c�xd��Md�+�:h����-��@T�B/��SЈbDA����6Q:(#��̨�(d�x�ƹc!����U �:���L$Q�ҝ��T�1�����A��N�D����L͚ր����0�5M�Y-�dA��D�sf�T9��V�v��cpU�L��v��!�%��[��)�$����A!���@��p��IdY�eOe�ݙ��O�\�F�% �k���"
Q�,�{�DT�Nx$Dv���Eb`���%(�����pid��`���(D�hrP`KЃ2L��t5�\��Qv�������7�؁<��cA �5�+Zu.�ư������w� �R�]�u7�����P��~��UU�u7�#��e;TH�3=5	]Sa��(�&��<^ܹ��/B���3��O��ͩͮ������B�n��BĢd�ksX�"
���(�s��T�3ȳm��	T%(�D:m�2S9��V�U�E��D�����sWl����dRX�|9V�X�.Z�����b�r.���s��Q��eZSr����	�ر���Ѽ��U+�c���������8������X��?GϩA6t�; �7�n5��^K�?O~�P���dD磹%�+�"b� �!V)�Y\x���6"���+�d�`�S�c<�]�16:�k�HE�����I��֖&Δ���v��B�Pď�{���ў��A��(m�cu0��n!	5J
�~�����Emc�l���W��qCɌ���Q*x���ˠ�9
�9<���)�C�� /*�"ȋ	9�ľ=X�r.�x#T��iY5��u��~��?����G�:����=���d_k�Ql?ҏ�w�0 ɒ��(!!zX1o�w$�S7S�,�R�\,���̫�$i6I�,�;$V�����V%�
 �-�J���Ε`@�*sq�9�q 3,N���
@�`P������54=�����W	A�!��a�A;��်C�H)?I�[    IDAT:\�!Xp�G�\dkK ��s�;6��"�Q�a�~%@�D�z���˗��;Q�h������c�zѲ>Yz��ׁϟ"��QSfZ�&1N�# d����.�paB�d�Ѫ|zuK�)5���d�778c�_@���l���Bi��>�����C�RA�`������� �}Me�X�B�^j��ߊ�l��ޝ�SF@Sp���3�)�����I�hoA!�g��m\�NN&Y�D����$���M�~?21���	l��beW��o����#p$���)HR$�$w�P4"&FG�A�X�Gs���l+4$�F�LtA�t���ݠ��0
p��JG�� B�A��+�/ekݗ^zG���ھ(]bɒ%hkm�u$����t���`/wHt-���E"q>O����N�t���Ô� ���$|�#���,O�"�2fp!S���ϩJ�� N�A`�#, n�&d�WLH�E�?��HO������ŋ���b�jvT����775��:�ʰw*��y-K�?O]ޕ�9v;p�(��2\I�7n�3���HC�cP�$�� I��C6�2jb*��8>|�
,�����>��06\t5Z笂𳅪 5zēPB.�EPõ�4��8��/>ŀx2UD�Q$zg�1�{O���1lZ�	7\�fk�Wǵ:��#���E�?:r���)G`硃��-�x����ã;�#����Uv-,��Du�+&�
@�T��p,�a3��l\��$P&zYyz��g��[B��C�y�wâ
��c}� ��TV�Y�tX@i�%@�v�D��U@Y��-�4�qV*W����0�\	�c�(hZ�W��M��6����bC�)��:"���P�,#�M�H�{Uc�S�rZu��]�	��3�o�Z)�@}�W>��Rp���p�ʁs��G6Th4���8��}��o>��aؿ��~���?��V�IB4/����FLN��,�)`҂`�jx�e,�衔�sO<�۞���~1M�c�馛�*D��g���7�#��\PS ���$w��^DnP��1�&����F�'X�}�u�xe�>���y��.8P��'j�3�m��ѩ��"��N�#51��1؊(��/�Xq��J�ʔi#�6AS��B6�s�4tI�C6@�9�V��ڛc�k�uwqa�c�K���#}f��c����KY��D9���?HC�
G�Y" A�P��9"�Z�p�U�#Q�Y����S?��[���\���Wu6<�eꛏ7|���d�i�҂@$ MsÃ�	TJ�W�)��@1;�s׭�E�73ް�\ȓ��$yhjld��H,��Iv�#[mꌑE0�[63����g^@�P������[�H	d�@j2-V�:{�m�$����՛;p����38[��,]{��W@r�'eئ�A��D��������y������yS��Tk�C/�:���	\r�%�l�z�vktVǵ:��#����?8pշ�9G`ϱ�^�v�P��S-ވ����]'1Q0�*�T.�o"��%�#��l�R�R�Q�
�\ l�K��rT(B�m'�9�@�E�Ȋ�\�^������4�4*�+E95����WЊ�4�ݧh�D�
�1>���-K�ߊ�T:��LeN�V`�~P����C�%J����2L�U��bX��L�?��+Ա@,9�C��P 7&$���-��L$��%�*��m���g�X��<x?��&*�}�4`��t���Lk |0��D]�ײ�*=����Q�5^զ�12
�5��d��π�l�X*@��	<��O������.D5�|7�|36c(�sL]���E6��"������T�E�T�RaY�LPW�;Zd'�x��z�����Sލ7��� �)@Q��U�j�J�,��g��Ȟ�"���U�y.;$�aMu�X�o�<�<�� d*j��D]'
m��$2�Mk?* ��	4�D$ B�}�N�8拮u�A�i�]�x|��E@���l�KF�'Q�i[�%��+��}���ĵq�X�l��kkp����A$�Dy"���	��;k�	t��E־׷�%��r�f-
~�g��l���PΎb�҅X:.j	\p�$j��^,�H2S�h�c�8
F����ki|0�0 �qx��[1�L���'F�}�I-�5 D$�'	ڃ�wd���2�vx�U��;�5�^�+��AB�P�3XH����,(W�4=�v�P� �v��1Ȓ��㞾1ZeD��u����^�I��˯�e篃WNc�*�{sVգ�C�@��!F��g�:���[�Z���O�<�'��b����
/ׄS*A&��$��<	��DO���p�t�qP���ȠU7v��P�FH��똶�U* �����#� ?'�(GD'���Xb�*�|�	m}:��lڜ��%�Jf��r�ʗ�YH�a�ݗJ�
<=�ʛE�m���ɺ� �a�����#f�)&��b��p�$���Vv%���*+ȕ�i��-�y���ܨt0*��}�0� :�t�Xy�ovF~ؘ��o����A��7�%΄�s!�l�g�����2,��H�B����e��6�\��Ɨ����q��^t�l���a\q�圳144��fMu���Ӽ=����b֬.n�p0`>�L*�]Z'J�2�Ů�{��w�	�=g_�_��.��
HJ��������]���2�)s�I]9��Ip��b����zTk%���E�SO�.*��ۓ���$ *�q9�4L��s��� �ƌǻ�5)���J����χ��U�YY޻��.��*�ou�< fv ��a��gwq�΁��e1Z��� �Z�r��]�˛,�U�އ�g����"���`�R��s�deed����^�w��FM�0�auLjۡh,��H�$��-�zp��I!�g�=�汒2G�J�r۝��ۅ�rx�O�����/���pR@��O�i�b���\S�<�{ �8a���F����s~<aC�]X�SĚ�ø��h���'���h��R+5S�.��b�[�X�f'~���J��W�F5��g^E����A�ހc2C(@�X���m�z<��w`(�̩Wad��џ�Eh֍6�o�7�o�V�/ƾ_��sN�<����@���~�3���
ȿtu���g�0�0��gc������oG�>���uƾͧ��ro�� ������?�g._��+�H3Z9���
 ���p#��9�h4�Q]ԀB�@�Ȋ^�
Zl���"Q��ֲm.���~��(���^\w^㤳��vj��T��E<����a������?[���
��3�x�)  ����n�4�2��ʦ��,����Q��"�`��b�m�q���.\����ɳg00�
�/^ĊM��2�-��L���P-���.�4iE	�Iނd
q=Kn�[y�A�t���.p_[G�M"F�Kk��ڛ��Œ�B�"�Ӓ֐�U�)�0�MZ5>>�n]��~��%��4�~�E�f��~�w�~�z�b�|.c�ŸE�&����j����b��G5���@7L<��ؽg/��z�7lE��S����ןy
�B/J��L�X-�6�hl݇����o¶H�r�y�X�
� ���I�.ᙢ������A6e�VZ�ۨ �I82ӖL$8�k

�H�iZ�x1HQ�m��^���_ܟR)G&$�t������kW�
� ��k4=Y''�U��x#Y6x�a8� �b����������1��a�,,9a�kXg�,�	�N�9pB��& s�DMp]L�.��
�M�֯�__B�4�jE?֬Y�R����"�t34!�2Ϲ%����|�5H-��Ncq~����WT��ab�����p�]��9�6��� `���ڮ ;Sxם�%\����쿁Q��с��#x/( �tk�)�q�������c�s��~
Qzjz��>^<vn��{�»�������tj�o���7�Hz:���@g�8y�B\��6"�-4bO�p_84���2p��KJ�N"z	@TGV&̪`4]���A�r�=��
~ri���8!`��=\�H$�MHѤ�^�y2 �,��y*H_iw�)fn��4s:¿��{����#����!b�éK"�g���;��/bX�e;�M�#�]D}lk�C4!c�c����:$�a�a�)e�F���m0�N��:�~��wMC����>�Z]�5aUy�����c<���2uɀ0��~cRH3��`����m��`k�L@��q���p��	���Ў�xշb@�[��ET*%EG3 ��|��p�$��%���f����|���mߎf������O��B���mL�v����6����Z�m�e�О��bSBt��	����~�d)�D����w%ٛ�.�������=�h���%��C�dD�BJ��`?]��$%)�J�x���q�����u�t�7=�TV��'%ڍ����1�^�\��g�O�����"lT�bh�t@�thS�@ދ�K#Ƀ*c�@"�T�(�y�*MP�y��q����><��;�0}M���ż����H�m�9�2)T˕D{����zN6�t6�r���[�)�qa�$�Plؘ���k`fK��C��-C��pLq��1c��4�B�^�<v;֯H���W���!�o�fo|��J���W!Q�@�^��S'��U�� ]�<Z�JT�<��,N�-����4�߶|� ���i��~M;�Cg����<���u��-�GO� "�h�- �+���o_:��Kb3���|v��)WtRi$-9�k!���I ��
��܁D�A �:ǉ��4��e.��8�21ѥ��I�҉����ҥkNp�Qe1�Wc�hH�3���NJ(�T�bn�;�|S�L
Z�FL��2��}d�Y�t�w��^��O}I
w=�2������>��to���܌T߀r	d������/�o@�!�U�u���:�:(��RXr�e���I�)��ej"�f��ö�W�ѨU�:&\f`0�&����� ��anbcWe���o���2�b�d�	4ԛ5q�c��Y�N\X�,��%�hb���N	Ug���BKb��k���LV�!3Oh�k�2Ica*�<ը�VДC�8fZ��+S"q8cw_e�Ӫ���l�R���,=�E��r�!Y5r%&�I��9��$`۶mزy� *
�����yYNA8X�r6l� 9!��)S�z��D�А��Q��6Yi@�5�q�N�108�V�cݦ���SO����p��$'�E�P���=	 T2R�x����ZV�eZ�� $V�,#��ߟǶ��x쁻5���
R������LӤ�esȦ2r��rI ����������0��'��M۶�F����Vm��RM��C�ho�-s�iu�^���bE�Ý�W��[6 h΢{�w?�hN���8y264a���}�FN���$V����Q,V��aT�"*Z�j&�]���bC&��߼?�}�#X��Go�L@ޒ�@砾#+� ߑe�l�Ͳ'Ύ�b�r�J�����3���q�ĩ;�t��$��8�K���ur�A�Z;	e�i��J;��:7�c�rAt aQ�PY�7�LL��#�Sy,����r�E��	 E�,t�ga�%ţ��r�"*y�i�k�U�sjA��b~���سc'�R���_��Ж��	lٺ�G,bZ:�ԗJ�t��T��"��+��.W��~S �LP�������I[ľ,\o��a$%�P��Dg"�d��i!�Ue2���KR�f[�I�݄��:<|������wAꈽ&�8q���Z׮]Q�S�
V,����g�$��ƋNH#J�y&&'����7�N*O��k��:6�ta%"́Oa2�))���'f�^���ݲZw�y�|0՛���7��?��X�P�Xl:�^X��nX�]�5�MS@� Y���!���'۷o�vNm5��⋘��R6�>�U�4V	�]]�BѺ뮻p��%����s%��0��x&���}��z��&E?�r�z�j��^Y
��w��x*��x�mN�6�"�*�����$8�	Z[��#�
;�m������@W����5���av~Q@#S�I��ض��	��nc��C��+v���M0���o�������W��µi��܆�z�JÓL������&�nx�ʮ�ɡ�v��+��y���8�Ȼ1��fh���6�:w9��
�ؓ{��"t���s��+ter2��teU߄� �a�b�Ҝ���
j�}�{�|��",]��7o��Po���~��V�s��NIg���+02:/T�ҕ��@s��ܳG��/��tM��1(��d!4R �{Ή�N,���b]es���C�RJ������pl!V�R K��2@Q8CM<H��z��O9Y'�L,�ɔ�?�F�'m!E�%N/̀������J�Й���d�0-a�E6��+��6n���k�ʳ��^��sץhX��)|g��B`U����.�x�E�p�&�z@!�)�f���;׻c�������u���$�0�hQ�ˢ�t�(��5k11:��k��I�.��"��Ʀ�����֯}G�G�-�����&��d@�)ҋ�o�Nx��JA��EI��$e�$������%,�+\���E�RA@���E�epJ^��v��@��D>�B1�A_OV�f}*������B�r���Ȧ����G�cdGj���h���l�S4ZD�<56�d� ��O�7R�v��)���gN��.iVt��c�M
(��{����>���.�KX�'��2�E3$H��!ŉ����3Y������6�5�i���+�7~��o�d��UТ6�@�EoO������S�a�}O��\w�	�>p/�mB>cݎ��ndgΝE��(n_}��ذnΟ=���u�\Ӽ�����^���)��?�ԟax�&<������ػ�=y�K�|�G:L�R`�Nn�F)[�p_E��-�l�u-����|�{�j�#o�����h��*�4[h�.rY��q�<v�T�G�a�"N�u�������Sז0�;#���߱z�v��sO�������l�ͽo�7�7�)���?�
��t%^������C���#����x)D��$�Z��!'M*�ғSE�aW݂��I-'W^'*J�����G���j%SEeY�(s�ҦI��N�Hlc����>V���y���v��p'��1ۄ�W9
J�6�i	+M���S�$)�8[��P"rR�tZ@F;U['N�����6���mR��hA�'wu6��ƣ�gy=�J	������ ���q�7NX� F�PୂU_�<��:+Y�{��8�f._��LJέbq��%��X�п��~{�oD�]�jK�(-UPm�q��)9�eX(�h��y)����	���UCC����y�߸_|�iY�:�8-z��z�%�ߜF�0%0��'�EO!��Q-�cnf\D�B�"�͎�0t
E�\��������Z,--��18��B(S��\�����Aל��Կl۲CCCX\���ÇUZ:�{�;�!oG^��u�V�ݻ������e�!�N?��l��K.���̴\���!*��bX|�X&$]��B��>P������2���,���8ACU��4=e(A�K�7iiiCC!m���[��w?�=;7�k��7rL~�3�Q�,��M�U.09>����	�i��@x�����SO>�%Ѭ<��+(�c�M������ܒ�/e:4�`J��e3�E�|u�tu�豪�s[/�0?7�����=�ah��ϒwn�ll�t �$��Lʂ��0~�e�N����9�Z
����D���)g�-�޲���<v�x���l��`g�O�q�y��
t �[�w��GN��^��T���j@�OUjb�M�p�"H�#��x�3� �3��]d�L�m�J4.1� �$_�����Cƈ�z[�Au���Q<��)"��]l�F��f�F81!��]�K�8���H���`�Cq��A(�}�m�a�[,�J���$�fqbpd*ᮢ���$�u�g��pB�tqR����s    IDATf�k�����,
 !���`-g<$ӣ��	�R9�|��n^q��!H��D\���7����(OM��S���!Z֦h���۟��ݴ�)I/WkR�֛��'Q+��m����|@�K,�X�C:�������$�ѱ��ħ>M�1�XB׊�Bʵ@�\
��Sٲa�zPL[8x�~�&��D�YǥKWp��!\�t���رcz�d���U�.D
�K/���� ����"�2ɜ&4�e���c�� ��ɦ���vx5������^�k���)�!*Ȑ���v��Z�:�l��j`HY��分&��bm̵#p0L[�)�-b��*�M��`xxH ���l�B7FG��̙s��lԛ!$^PnR(tA��HJ$��>��G1cc������Ө����X4&&&�t�,�K�b��^l�y��r�qB���+����H�g>�yĚ���y����>�����* İ҈�V@�6�!��S�V�=2�v�4����Eyv�SSx�G~kw=���ܟ�8�-����<f����K9yH���|��u�=�(��(�] N�U1��D`0�>;������=��ޘƁ[������i�yvg����<�+��׭��'T!�뺓�K �WN\�ɫ�cK������H�� �"�^��-)�/��2`�����+�V�Q ]]�P�BU��fҁU��u�i��$'C�����{�X�|�5�U [@��0�lK����hT��N��AP��-�C�Fco&��c��יo�TB��(R� .D,���ߕT�w]�m���9ڀ�MM㾶�ߌ�u���p\�n��/^AF*���|ب��[p��q4��<�����n6m��!p�رy�{��}[��s/��zK��K�Lg��"q(�ĉ��M���h�k;&V��˴��5ҝH���/�2�,�ؽ�n��.abz	�K�id�>��w`�ڵ(��~�#��^�����z�)�LNa�ڵx�;�}$ %�`���簴��s��	pbq�sBG+Ұ��DQ�ڮc�Y��(��8B'�Tc��-�<�*N���L�RȤs2���^_>����^��l�-���5���y���u���Տ�by����y|��m	��rU2P>��/�W��v�7d�D[ma=ҙN,�	y�T�:�ߘ)��B
�ޏ_�w��S���`^O�*)�~�J��z�.��u�/:`�6�=E5A����
B+v�$bll���S2����O�����(^x�$B�^�L��Mz�,6iha�E}v�z��"�:�]���7݌��+������/�]�-�0��-N�BW/�����������^T�n�G�8y���eT|-�D6���x����;���q�͝ �N�Y�ou�6oB��u�����_�)�$��pR�_>r/]�ǩkh�&M��;�N5Xh�~#	4S��tR��b��+Cf"P�!��e�o�G��d���MFJ��8�P�%V����	+II�� �K%�k��h��og�50��e�Dg!���;"����
��O�4R�˯� f��;��sR@�Aꖀ�7j=�n\��;;�׻%}��lY@~���C& �'Lhg2��,�8^���+v�ω�z����ۈ�U+ػc+�}��x��IQI�+�A~,=�����G��7�g�
핣Gbҭ���2)W�hTk(�T�9�ޤM�Q�גB���� Q�,�9`b��Ї�׿�5�=�.^�µ�y48�H���|�z�]��Gޏ�w�hz�đ�駟���f��ڴin��o�l��_����ɓR@ө�������ŵ2P���u�u�@0A��e��uvFf�'��k��r
s�yddD
q�uEv*��%vJ��H�"u,��s� �lٌ-[���b����e�Lͭ���o8�ѩ��?����_y� F��T��DZly�K�C��hVL��/:�UEܳ�f������U�2�P3���tn�(��Ҧ��M�e���PPN��+���G���}�+_���^>z#Ǳf�m(�[�4|�A�N+G:�.�u����9�V+�:���{�l�G��PkT��λ���o�o�w��ܥ8�b�}��<�z�b�<=z	����^t��y���a޷�g�pj��su̔Cz
������l���݋'�؊TX�] �V�l:��Z� �-tg3o��86O��KQ���pu_>t
G��pf|	UWG��!BX�?`���A�LAXQ� NCH�R�	vO҃^G�J��V��I�k��Ƈ�����Z,�8iPBXΉ���<���AL@�PD�4Dpl	����kR�I�W��� �et� �e��u�p�q�騭��a��Ky�2�,Ѵ�t���~ ??��$Ɍ���hO@��r���\���L���� �7���@L�Vׁ G@��]c`Yn��=۶	 		@t���Nf
 �n���]���w?���<��14�R
�J�&��6�!ԡ��D������ir�,V�X!� ںR+p������h��=�tm.O������#�?��K#�� ?�����v�p�F��G�]��\�Z�!)�k֭���:u�LL�A�������P�LB�Z��	��p�ͦ��ʋ�}��a�f�!�R��31�h<Z� �eW�D/�IC5s��LO|��_��_�������G���xnvIt �7�~�#F6�Ɔ��:�������ٳ(7��71_� ##�u�˵m�5ћP�͉%iXt��~��b����|=��V �- !0'0UF<.E�$��j`ꕚ�H�V��V圿��;~�����������)�O�
2i_Md��{�`,��+6Dw�L���b��F;�u���R�Dyi���Yh��}�<u4&-�,f�?s��rUj.F.M�m9�n���|8�ٚ�jh�L她�OYЛU|��xd� ���q�zs|�w�� �F<+�}������b<>5�2���gN����FU��j�B��J@�� NE��,с��T��',hTx��)�NB�,S������u��v$��mi�X�~����Fa.�9����B�PgGԐ���IQ�$��س:��"U	�3��8����^ϩ�>�<93�4'��$�#�l%��ܪ��:��rT:;�,���0��ο y}��|��C�o
@t�bжfG����}��*vmވ3G�#�T@��n��\3a��}�ٱn߃���ưu�&�\��O �sS�g�r'4�)�J��M\�Z0)\�dd�*�<?@Ww?�޺�=�)ix���c�8u�"��-衏�/����+��~��p��c��׿�\b��KG��� [�ߘq�ʵ�ȑC����,v�؆�~���THH`@�Z��y�$��={v�ԣV�,���剋�
�*����k����[���SN�����r`9^��������G�G=뺁_|#�/�!��Z���|���|������:~Ku�35�.6;'NX�RJC������y (գ&6�]���^�ؼG^���Ӹ���1�j���b��`B�a�� ��F�|V�?�b9�r��R�,yAj|�Ы8~���=���2������k��^���A�IO��C��4NpZH�5�a=v}�Vt�ط{�܆��O��{���|K�W�GbDd3���L�����8w��h��&vm���Z�(��g��_���M�xzKM!<o��|Ɔ�������C��",�[;��ڇug�o�xK����N� ��+pat:�^X���G������Փc87Y�9�bvy���v�I}"�6�����G?5"1�"� ��%�ᡷ'/�&`j�a�$�N�D$z���닸�I�$�t�a��D�5���@�t��p��L-jMJ�+�� �!5��<57 �d"��ľJ([�iS@����3�DB�gW8���#H[��,�O:��S�W��w<�o5��?�$ٞ���j�R��Y��-�p����J�G�e�g��&t����1�[݇;oކ��V��8�Ճ��0���}_���ղdD�J�^�~�n�Z�u:89�7]T�ٱ�Z������J1�{ﻰT��05��m6�����ǡ�.��)<��}BK�b�V.H.�����s���C�@�v�܉u�n�k�?{.>s�����ظi=n�y~�~]]="(oO��ڏ6 !���ߵki]����q;L{���0MIޠ���*`P�9>��5*��������X(v�����p�΃rLW'��_��s�:.���7�x��CC���籲_ea����B|���>�f�X������'����S��05]����~jش~�֮�ڡ>�Q��Bo!�5C�%�c`�J���5��E@��d�a�F���blr�S�0tSl{��]Awo�W�ƫ�O�����xI�a�݆�������j�%&ĳ�[�`���2e.e��C��V�Ȣ'�?���wmB��ªbv��[vCs�z� ���Lf��HgM jaG_z~SY��.�qy�yz�*�p~���3.j�P�/�1ri������ݹK ȁ[;6������2+� o�S�9�o�
���Uр�|q*�g����×pq�!.XQ˔4pf�muEoAwq�R4#�����N5<��	=�h�(��,kW���� ei2�N�A9ݨ-PL+/h	�7<̗�X,70�P	!|��]P�⥶'��v��|��'�"҅t��-8��SLQ�؅V�H����
��N�G���"#I P;[CD�ɾpR"����3���[m �~���O
%�|O;ܮ�{ښ���9^��Om��~�1��|k�,?�h��N���Y�-;��̫�М���Id�1�L~"�t���A�+x����1�\F	�����s��
B���r���@��7ݴ[�
'&�pm|LԤ� I�y�����럋��ֱw�� ��8z�L'#k01��?�0}�EK�����6ٸxq$~��M�đ*�v�K�o�>�} y��c��|�I�Fmݶ���Wz��]&r	x�w���1�����-�Z�X0�4F۴��69n:Cq_������=y�Zr�"�����I߯�������^>���/�{<zqT����yM�u��\��xb�y?��?�z���H(X�Z+�K�i��D�t��ם�i�dD���_���ð�P�\Z.WK����I�6n�$�/�ZY�)N��6n܈T���S�p��Q��ĚrXՋl&���9ԛ��<��a���X�z(UB�[��)]��2���A&�E�^F6e�WΉ04� �4�35|���1wi�w���{���!�#=���^��z��¥��o� m0g���Ѫ-�KO?)BޏGN^ĵ�Zf"�� ��� W<\��bZ�%� ����x��w�]��A*\���w�4w��X� y���!|�V� d�R�8;�.|��9�ta�fk���[��PoZf�:�.�ä��h�RfJ�8L�.⠄������>�A_1�\ZC_w�jYٽ.<�����4�bX�;��n�Q�X�i���<*� cӋ���F��P,��Vo�-���ZJ:�D2,�C���̤��lh6�.^zS	�*��5��R(�9i$`���S" %g��[���
lON�EQ2�F�lZ��I�&ܘhh7B��yH�O��r�Bq�2�$Q^�e��$H�#:)�kz�no�䈩s*�M�4�5b��-I4�u�6�}�<R��*S��!p6g�0#�'��|J����W���V��ꕒ��Y��}�}�Mزs;���Jq�E�ۭ"��xqDܟ�|�)d294�M:5�]�_,	�/[��>��������1��+�.����?��AV�c�`/��66�_�M��t������*�{z����L
�o����x�dd�\<1>�����}�l޺?�/
�t�rN��X$��<���<��P��91�)SQ�"���t�T�d(�/��%8>���k����,L�������oٿ�Y��O�Q<?� ���W�J���������w�q�f�#?���ܥ1\�^D����L+��-�D�"�>��-I�&���;�M�ȑ�%<2�q��[���G�2G����{�m��m4̝>}����b�� _Dw� �~����J:�]���,�'��=-\��5h��%9Q�xo�@!�6`i�XϮ(��FsX�o��7�2{kWo�=�Gv������__�uC��Z(�a��.����J;�[b�0>��3X��.LV�#�0]��yxd�
eR�;g���>�����};��g��m{:5Է���Jo���<o��9ܿN����U4I��Lxz
ϼzO�����R��oj!6���l Ҍ�_�4*S#�-@oWk�
X��F
Mt
i�vl݄�}݊��p2���%!�S���A��@���3Ͻ�R��l�*ߝL���\9�|5��t5/B��z����L�W���Z�#�\�дX:)X����`P,K�5'Ig,���I9����8M�FSv�I��(A���H]5���O@x�"��ΐ�" �����Q�,�w��i��(��KN�r�RۥVC�B� �/��3�i��/�I�-����+�/q����޺��_��N��b��j�2Ŵ{�<t ��ܩ��6��cM�I�P��Ѩ7����]�F�+��m�*nڹn��W���P�X�R��@G;�`��Z�� ��0;݇�0�c	<3�r,��
���훇��Į��1v�V��A�@�X�2����2[��n��j��V�� �����}6~�k�b݆�X�i3~�g~�t^ָ�2!݈�y�pb�B �sGb� FI�e;��'�l�Eɒ%W��ʘ��d2���Z#����9��?��x||R�_SS3�?��?���"�^*�$��?��b��8*.>�xY��Ђ��I}�a|��8�[ֶx�zX����"���M���"
B���ѷj�y�9��e�ZǎÕ+WP���@��Y6R錸��z��\�ba���N&# 4�<�� �iM�f�P@�[�#�)�F���Ъ]���m�����t�D��0����{ӇV��|X|�]�K9{������r�c�EB��3��JӥW�]LVZ��d�H�%�*1�SH���,>�=��$	��[vwj�NQ�Y�oq:7Ϸ�p�?{k� H�m�0؋u�F/���?��a,x,~L�~�b�M�-��C�!j6�7Ly�Ǫ��sȧB��ؽy��B���h��-��k6�hT�l��<	B$_���#�d0�j-����J��+��x��8t�<����*0�P�ܒ���*���Ў���;K����[T���e���C��A�H�r�hl;m�� �o�*hw���������I��D�x�����%�6�KBq�aP�$�	��rNE$I[$������~^�#K{���vG^e�X�)�sa�k�a�Ţ�z��Ŷ��p���"B7u�N�L���ְ*l �K�2"T�ו��Rs�C6bŻi�n���eҨ,,	P��/aq~NV��
�Y��+V
U��$:�ı#�K,�u�sZB��4�(��ݷ�Pz~n۶lDOw^ �%��rX���rYlۼ��El۱�:�o�l8~�pL�w*�������p��죈�iIs������Z �h~�)�u�!<�a۶������o��C^_R������� L6
>���cӚ�t��{�%&��z3O�kE�<mnI�]�G������Ǚ����e��`���S�M�\�ޓ,�%�\��:����Ri-W�����`��A�q��[7��e�-������	��c'�03��U~
-�M5��M� �+J�ݿ\���&�]�q*�36 8y!xW<��8�����b���q	+�uܺuv�Ei|n?��?��u�Ȁf���ҫ�q�5���I� &Z����"��z�Z�<�f�A=�!׷��Ǒ3W0��bL�@�0�EY鷈��CwD�4���0��x�{;5�q.��    IDAT[���w`:7�w`�;�x����q�����!038ta��#�V��E�6�j��lс���=�n��N�'�����U�Vw�w���5Z9�*�FW��y	,�lg��s;؆=6`j&��}�^8}�B��c�}��qj�*F��7�5���R�se�@��k��rRN>�&�����6q��7�Ē�+5ih̓�@j_t�J H�'I]gy��TbWz]�OU;?QtTs$�L=&45�p�=�d�ѦP��F�gUH,�%c� %�' Da"���Ӷ.�ζWu�a�階��J�&���t�8��Ķukq��!�� �$��f-�,]����x�k%h�J��4,����A�����"Vnߊ�N�W�uq([74�ى	L�^A&��/fi3��R�M@���B7͖����K�vpS3ahp���V��zE7,��U+���)~-,���z�*�~�>��ٳ�q��{�'�]����S�O����2y����#G`3��W!{B����0���*
��C>���Cѯ !(% �@Lq#�T����A*�k�@B�>�����lx�7�C��D^w�lCR��]�W%�����ħp��B=7օʘ�Y� �f�Z�؈�y=�˨(a�a�WV̎�ـ�I!|�'�~q�1�|��.hV�.p���]8��!�Z��T�n�vy���l'\��MG�[����f�^�/e"!�E�f�w�����q�!g��as,j�{�&��B�9�M����[o�ݻ-׀Qx�[�V��7��������4�wq����=pr�����Hu��n��t�œϼ�zh��ƨ|��h��9��F���1M��EI���0�x����������7�
t ��t�绺�G.��r&jY<-�gO^�߾r�s0l: �'���X�}�Y���ż���]�̓:6�pˎuؽi5Һ���`��Q�ESa�U���jHWܴm��В����.�K�uua뎝شm��o^8�*����:]���G�7�T�0[P�kb/��iZ$����p����C���9d�YZ�!"C��'.ZR�K�O��x�^j�Y�h�a�V��U����ۍ�qɏ��p( �%Y��`��^�ѡ�PX`�(  i�u,��h��U �ڮ��8���n]M���Ir}Hj��)�,�I�K�����@بb��8��h5�)T#�RE�p��3��J��r	`H8�*bxM��� ��͛�4/�l���;Q������ؖh
X�g3i�k5��F2A�y�)S)��M����k����[vbx���G0?3-4.^{�zSVB���kѨ�$�cppP�����)�:v]��P�2�,r��łhTh�+4)	�z[]5�)�_��s�6`�
O��\;
�(l�Ћb�	B�j1!�f^�rK�w���R�G��ɉi�*UYs��Y�������J	�p��n
���Z�G�g ~�#� @�T� ',��_��(:�G`BZ#3K��	2�`�ON;��S�ajv��Ⱦ�]5��/��`�"4q��cɖ�C%˫�� ��?� g��$�/�6�t�#������-�����T�n��`�\lYӍ�9��L7mĎ���^�# $?�Zf��>(U/�a���n �O�����i�O�bbbBht�Zg.^�l�C�w-�����J\���k/E�;�Z\R1m[h��W����Aʶ��e���x��a��x����^��wV�M�o�7�7�zvv�M���_�O��� ��+��Ա˸��ނ��h���k1,�Q�%)�fy=�pWll[c��{�s�Fxӣ��_�l��j��dvC�QGੂ�bT���;SK7�S.T C�j|jR����<���fFlG��O?�c���B�i`���\)��l���-S�IO�LC�,�
PuOMC���`�+G����BBA�HW�]Yf}(��A��IQ��W�(��\7�N(��B%9KD"W]q�w�ƄYZD�[�ʄ"Hm �',f��AR)�X^�^WS�#՝��VlэI����s�|�]�j�y�F�|�Y�
� e"���>�V2	cz����I�����k��5���+�ۃ�]�4LĞ��[�������ǔF�01g�,�V���y��'�}��`&��"�8��������4�vg�s�l޸'����Ź���h���x��~�#��$��p��e���˘����M�3)M�|^��rRp]7��D��U�@=����e�0�]P�>9���E���Q#�b����G8�C�Yĺ�˗/KB��d =���a8�� ���5A�����O�!&�כ>�4+?6P�C���iH@�H ڂy�M�����H	�����?� `�h�� Ȧ���E�{M���U+�s�V<��/�ymJ��&�%M��
������0D*�U͊d2�;��: 7KA�$���5QR,<6�I�F���l��nظf ����1��]�mY�9�7c��[v���}�}�����8������o�Y����e��͡���B�%�Nc�3�X�E�B�U@�s�i31�$t�f�u��D�`v�Oe� �F� �Y����ݵ騌�:6�o�O���7W����\�ζ�~+p���������;Nu�ˇ��d��?�-uZ:4&z��3&����;֣��cM��Ҏ�o�C���[:Ҧ���^�!5�G���:l�DB���FK�'�f�����ی�ջk7o��]��?�>��g�?�
"��-G(5L��,�+��-Jq�u���ܼ��u�P�I���s]�NNJ>��Q��i7�=eJ�D@ nXmz�$����)H��!Z�i%�H�!�F5Jl�u6���[Kj�:��4"	Ѫ��X��,��=礅�����M�a;¹gN���rC#@e�rR=mV�ټh("��b
��i��^{�n�I�,-�����J�B�|�e'�R���Ҙk��ΦA�e�Bq�0jf��4,�Dvmނ���{U��&��<\C:�!C%���/@�s�0���s��}�I�5k�[э��<���H�^~�yD��HR����K���F�*��w~�?��_���4Ҷ�cG�`z|�lV���.�����g�-.k�(J��XҾ����J>�=
�!�kA0�1h'|��f�����6Z�8`5� ���111�r�C�2D7AA�5�\F(lk֬�����L^���¢�ݼFt� a�R�5+kLJ'0���LPZ^�l��:N0�N���&c>�,d�{&N`}�=�m�^|��O�:>#�!m�N�%�n��;�W[�/n\ˮo�ۃ�p��Ѣ�"7� $�{A7l��@&堘M����vh�����C���`�^4�(����{1�z=��35=l��Ç��������� ڕW�-�����]��"<�3�u�-��lx�$��,���%z2j�-�u�}�>ܺ)-4+x�C���;� ��q�޵���W&t��۴���۴���yk����#"Bg����Z�|n�~�U\Y� ��X>E��އ�9�9�,�X�gcC���ޱ�m���qL�����UdL=ŬP�X@
=(7�5�b�ʎ1�@��J׍N���N;2i��B��$��u� /��	I�S����wⓟ�>�����Aa`#FF0[�19�a~貣gZL('���9J�:Lh��tZįf:#�!����9�=�׮ېRL�[D��ƢA��p�T���8YpI�c@�R����E
�n����Ԛp�)X�-]�Tql���G-�)9'�e#e6�cR|"hfԧR�q�"!�-(�֭��xyaSSH����:'b��m�q��+h��`:9��5ju(�&R�8�{��-�MM)�Ո�t��kP#+���^ �m{��:��㯼4I���,s�4(l���؏`:~�d����"�Q�Aqw�D���t�j���kW��M�Y�8�Q�b	%I#1�� �&�e���]���+h�+�ǌ�H1H�9jBd(��Hwj��6MhY�L����"����!Ҝ� ��0�+Bww���R)5�	�{�^���"��:R��KG6�A�m
x����b���Z����q2���U
�)�O�x.Lw�*��<'~~�Uy=��pe(�BP�B�LVWF6�RӪB>�;nه���<�όȵJ�H���|p;JCCP�����+]
��X(sRȜ�cj@ a-&���F��u%�|?I�Mt�m��:��,z�&��)bۆ>
H���;������ݿZ�Z�U/š䱸HY..�9&����Iq/�ꘚ-cz!����B�w0_�qyj	sK�P�^�ZgH�)j���\hž�i޷��A���{�.<q�nt�.�����5>�;G�VY� y����q|[V����q�w�p�𙵁,�L�/�9�kea�)�B�p�9����z� �]1���a�`�{��ީ����Sq�f<`$��L���id�T����[X��G��������u4�-e����n��5�SP�ޞA��(WK�]\»�G�|����I?��/.b�a`��]/�ӭLA���
`a)�!�����&��XG:�g�9�~�"��]_
~z�׫�tw'	�:��u���TN&պ�L� /��m'�z�F��`���fǙ CD�R�k���c��U1b��*�Bͼ�H��Fw1�I
�.;�L�4�ɜi��pJ@�'�*@Iw��֛Q�fqq�"h�J �iT&��cƸ����x�$ξ�
`��5���u�4Z�*���>r�Nhl�ejap�o�u�5��u��������2mM����:���R���r����f9^�q ��Vy*���0�F��pO=SK&MN:Mo�9I�uɹ�ΥQ//������ W�X�9�����d_�1�'YB��%Ӿ���'����MS �\k4GN�+mJ��?�u)Λ�=���m;0=��R�)nЂ�ʊ8\ܫr٤x'�N#�d��ò�h���F &�G��z�SCK]�湓y	��N?x�����*�T�t�}x]�2 5��<�sP)����G߅��}Ǟ�	�j����xA�5��&�W7�.��;G�B�le2�;F�;1p ����;i��1, P*�e �NK�E�����2�m�rطk-Bw	^����lٶ{�:��]���h����/����8�bV�	��q��o��Ě]���,,;�0����%,T#xqf~B��(���:�\���R�SW-�RNz���]P(����V��'P�AW>;j�=ލ��mAAwq߭�;5Է哷�"o���<oǳ�9�o��/\���Z�*�����Kg���a�� �3��2�61�:�l7o.��=x��;��+����x�+O#c21`gS75)�#�1�P����"� �ֻ,�}7�Pv�K���ǕK��ߝG6�I�X.�l���7Q����
������!~�w�O?�*Vo�%��l%�B%��b�Єig��#�ΤpH� ��3�FDKPj�M��S��2uTKK���a�`n޽+VI�K�D�S�[�{��]������=��fM����]�Ь��U(
�ūפ@�>W(�'8�x;�e,��}dQ��DL5�q,x�8,�Mu/�����ly�eQ�]h���N�H{�F`��\%�䱣��-���*e�k%8p ��8��1 �����߉�<U�f�=�Qy$� ���Z[�,�T�}��#�.xa���[-�=q
��Y�:C�q�#�����q��	��t�ImS D@�ZD���V��P�d;X#�($8��dl��+K(���6@S![�Q)/bՊ^y-��Hۛ���Z�:%�a�|�bW�]nZ��І�9;�B��IMB���sJd���]��w��1�ʈ�*�5��Q����>d���v�f gGF�JwIQI���y�mKL���Ǿ(��(��%!��"EBA�iI�� ʤ��$�1\/R�1�Tv8�M��5`���ghl�u�z��p�}071�CϿ�ސuʝ �pp�A0��ے��D������3������h1�fM�nS#�\o5��P_�7�C�4�S�È#��COQ����К�x���ظ� wiVrp8�����\��+���O^,��2�����g��c�U.�̙S���A�R���M���Ĥ$�k�^����yT������*��O���J��~ %��"�\�)���^%�F5<hz�MH>��}x𖭰�<p��Nթ':+�-�@�����go�x����.�$�(๓W�WF�ԲQkFR��P�uaF>�h�ש����܆�z1q�8^�ʗ��$4ۄ�Ϣ�Ь�k�;0�]���އ�N|-~�#�8l��tg2X�? Y�S��f��g�>l��>̍��?��b��׋BA�.����}��kH�3;�� % �b��P�8�`1ee�H�:�fZ�!���'��C9l�iڨ'�
l�j�n _85�_ŧ��i8=+Q�Kh�.�,�-�kZ=hbh�*�^C*�=Յf�).�;�(�`:N�(��k���8���?��L��\��+u��<;��.K�$0�b(*zL��sDrTD�ĈA2,��9��ɝ��������y����������B����k�LO�[U����)�y�D�	#Ӈ���WD�U8l� �^�]=�b�v` �Hwf��٫�����n�'S�n�zlٱ�GFQ*y���;T���aYzJB&?y2(>����8�="͊�Z��p�lQ�š�[6�F�uШ�%���������~�Z�c#r�dؔ, ���ɵdH�x{d[_�&p��x�0�X�\X	z;l1�����Ȉ�����@�/��*�Di���(LJ�(]�λEyAN̒Զ!]���D�D�y�h��rIʈ��o�)�;��2I�j�%�� �D�f��Ν���׸(U=dsݨ6<�L
 H���JD�tJ ����Gd��՘Rҙ��B����
f/K6��k3D>I�������c��&pJ�c��$.3g�D��i\�<�t��X;MKo
���i��z%��M��QS�(�b�U�J	����u����B�ؚ��u�����tf] ,�YA��'b��g��L;('�?�3�����K�f7�K�)�w��ةj��$�|X�0��¾ٖ�Jq�R	��	�߿O
�I2Yn`�p[���L�M"�s�.
��|�@�a`�\G>_FKpD�f"4�����c(�����km����`�:����p�	���'q�	��v??�)��jj���zx��5�z���
�x�)�X�����J�5�pˊ�(��({l{��W��#��Kz��Ϝ�.s����8�e3f���U�ѓ�m���y�>f.Z�܂���gob�J�g�&�ݎ��0�z�r����*H$]�C+���W�
��A|����>4�,�A
#`˞	����P�D.RׅO�J&�2$e�բ'~�c���9l.��2�U{G��kH���e�v���1'.��o_{=n��	��ZܬD_rmի�y�t>��w��Rn�{����>4�΁�W�k���",ۂ���ՋP�"V��c�hu��.^���q�C+1Q��7��u.^}�R�B�ViI�h�#�MGF�"�@�.gW�0�y�
\��kQ�,�Ff�6^E�Y:ؐn�� m�B��h���Z18���,�}d��p���|����f(@�.�Q6����=[7�Q��u�@�Vd��1��W@�Jq(��.=u�@����LWV<�r1���Z�:ØёIJ��J�(?"h��+Q�dC]]]���iD�mb@AĄ��T��E�J�q�#E�.�&��-��1��!��6|�/-LL���v#�ٍ��c�p��[��y�q�
�B��Ň�Mt���,@�7(>g�B�f�`�*������M���*�ZpMH6@R�����t���藉����(`�Y�4�{�j���j����Ǯ`���
j�����d�f�Z*�Z,J�%n송w"�y���9�G�/��V�@2n����@Wn��Y@�/�n��    IDATUp±K�՝���?���Wǜ���?m::;���v"�逛�/��[|�����t����CD�̓5#�*5�z�"J�&'�06|@����t"-�i���#_k"��0�}0=����h����b�ƽ(���"H�=6d/��Q���X�5�i�&t��d�\�_���-�/9n	Z�!���c����ϣ�̩S�Z��y���y馾�����\��.@�$^��{pF<���4N�~UE��I�u�ڋ?m<����w!���Ӧ#?VBG�M�F�"(x%��ߛ�_ަ��غa5V��!d�6�d�ɘ�w7Wo؈S�x1�>�t��&���[�)X�uM��4�R�%R��Y��H�N%ĜI)OG�F�2���㉇��<�06W�jǱ|z���TS�K9�N��"���M[���^�I�
?����oo�K�����3��N+�'?p>>��#���-�޾���~�gx�����<X�E&'Ȑ&��Qt:!��Zx�f;��k��n~�)�L� ��B������b�l2������${Î��)���*57e��}���6֏T<����p;n���$���@"��xg��mH�h��Daɏ���QY�:$0L�V�T(1A��D:+��i8oyM)t-�Z��aԊ�������P�Ia9bLJv̰o����g�u��t��<ߓ$,��Q�*,2���VlL�G�N-~	�>�j=<ϔ>�X3锜�X<hȗc�l�t1�:Z�E��5��z��]9�b���y�lU�ב/�\}�;߃��f#����o����`9	1�ݔ��1��fe\vAC��s��h����M:"���%�0���K&4�h4�ܒ�rβNF�2��G�`r���ր���M8�1|���;��D����H�'Cp��)�{��`��8s"�D�A�c����C�����H���
�b�8���Z��vE�F~�߃�d���8X1����P�l҄��G	��#�f��Ɯ����_�W��9�SYtttHX �S�t�LZ�r���)�$��>�8��Z����I��5'3İ�L6+��b��1��G�Pȗa�)T�ۑ�A-La��o�Qb(7Z(�=�ʣ�4�xZ���S���3�����L7����AvO��0̠�7��4����a{�x�	S���0uN�=+0@�{�y��������*O�h�Zv'ݰO �P�GC��ΐ�ߤ��m�0;�pY��-������*��M�ն�8r�t��D�k �Oz�?���ש��0�|���X�;��J�)bXr�1��{�m�B��Ս���m�++���S������B1�R�c'S��鸴7�c�z<��[�-U�F.���N�17N�XW�U:n��������߯��>�XSS�������vةn��nT��0�?����"�^�k�&�2+���&�K��K!_�$n��M�T�"G?��5�U'��}7�,հ�3e�,������+~x�LF��K?{�;~�ώ�5o��X�{R����ȗ+����jȤ�8ci����T�/K����a�p���w�a�b�j�6�sXi7��|C�I��E�˫��H��W=VĈ�K��C�!��قΒʘ��Ӧa�ƍ����t���fBB�w9�,�J�##�ʉ��l �̄+�'ʡT��d"	f��Zj�z�;p��'��{����(�̚�}�v�RlY:�Y������� �H0�9�@��ȉ��|	\������b�l�h��f�̉�tlH7F鎴����Ux�;�)�/�qV>��}��`�I(��ER�?s_��F��f�A/�!���<��`vw"�ׇ	�<p3$�8�-Y��z�9g�F]"\i���Y��A���O?;&;�n���Я5F����}��/��n<��b<��e8S��.�����acl����7�Uݽsa2�Az{�}&1�"���J$([#��m4�*�:Rf��0���#��3��t�TB���4n��k��.�Hq�b$1� �v�?�k��Ɓ �ut9>�f,��̳�>@��NC:_�h�i�j��2(�&���h���I���Ã�S3>��v�E�h�a�-��d���tK�t�R����%�l���ڗ��c!V�KO� �$o�S��\��0�<��C�Z��i�lڠj~C� ������������!���*�F����w��/^��dk��R4W�H�s�4���DG�l�Z���/��<s~a��Wưk�zL���֡ݻ�ݑ��~T�Mt��Lfq��Ļaegc�d�}�-��_��!rbZזN�J��ӒØa&y�~�x�K_��g�*X>�_����\�����0�w��[{2q,_<��G��3֎��}Y㩚R���x�ՀՉl"�9W|�B�x�mlW�m ��@5f�S��y|5�D��������U�C3���o��R~������ܻV}� B@��ʟ�Lfk���+��s�d����I��n����PB쟘@3���2^���N«�y	�rI�3�ԫjQ"e��*u�7���zT��\lΗ��%Z�����:����$���r=�e���� C�r&��hY������MbC16CG&�Y�Ӱk�vL������^LX�-�mPp0b���,@"���,�P�=�0{`��!��
x��?�W��l|�[��_{��-���>ٱ�?�;̤-Ժ�B��P^#5���S�ZM��DHV@46z>�X�]���!��/;�, ��j�N;�4\x��0}��ݳ�����xo>�<�kd��0b�x��/Җ��;4����#����N}L�����.*<aE���w��-���{0��D3l�'[����	��"mHgX()��k�����m�w2��Ĉ�5��zy�4��A_��K�Q:�W��B�Zr�s����"LG����̔����C�עL4�D�Eٝ7��Ď�"�$��ꈫ:�[Uk�ЕI w�qmIMc�Hg6׉�/���}J�~�.a� �*�y�֚��(���5�(�<	�`pEˈ�\o!4�3��Z6��j�+&�R�)?#���&߄2\�*&�T���iu|F	��Ś����N�&�H����ac��~���#�p`�e���/�Y�-�ݘċ_0Մ�7��N}��
�������Z��
�޸^�M�M�0������oÎ�
��M�B@ �f�������G��~z�۶��d�9����C�̹�1w)f.>���5����NL��Ayb�֭A�qd'�o�Œ�N�{��q᧾�C%t�\�e��v0Yd��l-�\���f��fd�n���K���S��_�P؅�����詡�*�{�ZIX�<1�7�I���J�?؍w��\��e���W��n$3��n}
W~�g�´�����>�>�����ƺ����3�;�J���U��E߄�=�ЀW��-ij5�M���6q�MW�/`qo���ۮ>z�հH�
?�֗q��g��v��]�<�~�l'ʍ&L'�\��ã��f�p�t��m�����,��q���o\+7��]fT�W�R��.6wۥ���>�5#�9�AˍhD��'%~�ug�dX'�!�z.(��hY���c���ؾa3&������]0%ٌC(����O�%��4<�V�Nۙ�nW��T��׿'{,���p�o�]��o��]���+�n�*̜1C�`��h�=��e����i�I"�A� ���y�f4���η�d�>N�����ʕJ��qJ�He3�$S� �����Hʶ�~s��Ʊ���|���X��0��Kx�[�����d���Hf)q="36=�+�OiZ��S��:��_LGk�)#$��]+�዗�`�/���1Y���Fr^A�1Ӽ�L�"�3a8�\[���Ȩ5`Y���VL�H�$���=4 ��3�b��~���^aT-�}��2m$L� �{$�'��v���xoc�V���k"^#��D�1&iťs���ӑ�k6��5��<�UG��9�!;qSI D.E �"��dS�d��|��l��AP��X4�P��x��]�<T=_3]nRX�Q��A�"h3�hҗWj���'�5إd@>,�g����lȈW��.���=�C�pR�Y$2���_��ۋ��NI�C:�U���N?z,/����#��>�V`j��+0�����l�+��+��z@�\�Z(6\���܅�J�Fg�Yث!g����i���c��^b\}ɻT�g��@�v0�d?�D��=�<k��:U+���U��C���L"4���%i.;v�o}'�O�q�U�`�j�w���6�a��&&=4��D��	�L����iv~'1W_q1��;
�j9&���W����#�3�x��JMOJe8|q�P5�[>�s6~���K�+G�������L��������'.�����6>�D��L���0�t�=�?o�Ŧ�D�E�pJ��7�T���o�����o}B]u���8�R_��}x���=�y�z�ǿ��:�)Y�U(#�hgK��������s𾷿��2�����x�'���Y�a<�@�2hѯQ�T`���͚���a�.k��^�zH�	�@��;�Z��ͨY���2�W�%N����n�ٲ��1�ju�׍b���6b�]w͊h�A�'��u%�&�*��p�׿����Ao&��^�ѱ(�
�/a���h"r4�a_
��q�o�	~�<�g���,MԬM����_�ńaA�iѫ�hy���������a�]���A?�LKJݓ���F�	3�hp���5��8t/	�8��4z���x�i���8�$���y~4}3��kԢ ʌ4�d�t�&�Y�I��4�'�r-t��N�s)%cp%Td0B%�l��V �Q���Kr����{C'uIy���5	�bff�5L4�5,^0�����wa���Ţ�F83y�|G����5�i�f@w#B��%�#{\^b��$;�B�e$8�9-�4�<�0ӏ��5�ך4�S*h��#m?��e°�gj�R�BVR�u��P�{(��"�"K]�65c��2ŋ�����M�� I��(����#�\l���Tku��x�-�=�����={�n�z�����»�|N>l&,o/9q*�y<L��!^�C2�c�z��8d+�r�*UgZ�a�7Tǝ+���U{��%~���/�Ŀ���_v^���~��0�!����������Ö����h��[T�`��_�8���C�R@WgV�ա�<�}�ɘ��\��+��S0��(�-)�����a�5�i��N a�Í�4�^��bnR��*J}��G�o�vʔ!� �њC)ͨ�y�qĂI|��ߏ��:	��
���O����a�z`��Ջ�.�N�5��y�R����Z�gTUn��^��᧰�XE���J����7ྛ���3 䒟�I��Ϗ�a8�&'�}>��c�]�e5�/c�f�Z��K��������a��S���9���L
��}��aa�o�4���Z�1���@}�+��C'��M4�
��͡��0m�IC��&����A':IA� �'�X)lE�U��@�d)/�����R!�T�q�.
F5+B�Û��䠟�:N�����X'*	 �Vsb�C���HĀF���\^� �r��Z��kh�.	ٷI�A���mO�����@���j�t,�&ЩWR gQ�8�]]�����������M�F�d�Fs]�X�̞� �=�>r�'�y�DNҍoW�B;=���ؿ�������x\K�!�t.�:�BB�Y�p�N˲��o�q}��Di����p��L^�,�)bBB��� ��3��`�>zz62r��U��)10�]aԯ����bHs ��c�O�6�׾ۆ)^-Xji�	[�8�7dHW�0?�Z\3���յ���r]$�EV���%�S��� �9!��1�rJW:oBz�x�dd��@�ހ��Ĵ��5��q����!�5�?F*-��7���R�f���՝��O�C�0Ri�\��0r'���=r\,�7���Ů�v���q �|�+q���ycx��GL�P���xꅟ�+0��<߯�����V`Նu��ՠB�M�j����'�Ț��* bRF�:��'p�YGbQN�_�۔]?S͘��^�L[��C���mP�_}���.�~�>�K���$%�T�$I���w��0~���0Ѵ${�s�ǁI�V���#�F�;@\I~���_��^t~��w<��G}��˯�]+�����["M�?Ӊ(�����sQXE_gG-[�R��O�E�7`�S,�Ӌ�~��8�_ٟ��qϰZ:k�xp��n��.�t���,J1�ch��_~�,�� _��n��[��N��\|��ˍM{GԒ����ڤ>���Q�2�V�⃡�$uI��]q�`d�x�Wh��z�d��}�"��-��*�$;��@P������ Ζq��j��uG�^�v�&=�����m�d�n4�U�ʕi��[�9��#e9@E�&�oi�m[��%�	w�e�����Xh���|�r�	pU��W��=�R:��\.J�M�zV�v��J2|K�fF(�m�v_�>?}���B�����W� �g�"��r�z�5[�1m-���f���~4��Ȩn��>|዗��d�T\���86"v)l��42*�4XL�b Cd�o�\�Nm���	d�.�'>�!��{54��D�zD}����0>��C*��|�&�fĘ���i�J�����D�%W�� ��6�[ô0~�/�?I�j4�J5{� T����8vn�(�g�@��|U&t)I�"�Q����X�{����43'��dkMK�v2!�*��!�X�H�R�(
�r3�&�#;Mb!��@0!YY��,L�d�u��G)��YC~>':A�CJ
	��,2H �J	Я����:�tN惲Qa�؏�P��`��Alۼ7oC.�������
�` �:���r�!���_z����'\�����M�[���7�B�ѐ̯Ϡf8�k�j<��.a@�����0�3��x�ɋ0h���=����[l�D�y���]~H����5J�54�y�w��QϏ"��ѝ��R��m�8_����?a��}���cۈ��W�DEq�dLg����ҵ��ј�PۋW�qn��'��ډ@}�kW�G��L� 42�S� ;ߡ/�<�h0���C��"��B��Gv�I�z�|��Gw,��N���&�_����3��c5��J`��<.����9\E��☁��Ӫ��믂[�bnOZ���7�P߽�N�[&\���3����e^O�q���꽟�
�ψC�99��DL���%la�@��v��Ʀ��Z�K����}S���`$s(U2���k���i���,�.�����M�,&��E�����'$��;�Q	#�E&@��*h�w�9kq�Z���-ܖ�% ��G�r�4�b"+:��q�W.�Y�c;���/�={�4R��`��z���9�26b/D��jIB�ɝڠB֕ă�%����삽�N}��4f��p���f����I"Ao��j���p�/n�Ϳ���>4|���]�U��#�ǁ��F�VM��$�dB<9�#0�o���_J]Pܖn�N����HO��ڟ�gxiL:�03I�����:Pe�/ϟ�.� &0$���yP��~�o��]��'���1a�l	ER��q����NĮ�[���v8&�5ap����:.W�Eʻb&!���D`��g�VF	�����{;h"�X�f��z��e.K���3GY#���\�;��Nl(m��@����Z�F�$��E����&�0�{U'�����2z[7�Htt�����M�aiym�7�̙���ga���ضc� ��k 9zv7��>��L�ȡ{G�z�x��!����=udS+�_�M;v(Ʊ6�)r���8\�ylvM�шq�U��v�8��.��| ����z	6���]������C��U�϶`�������p��t
����$��p���    IDAT�����3k&*>Fk
+����?��%�Gh��,@�R�fM��!2�������W��cz5C����0 ��ڄ��+�����Հc��ʹ�0I;I�Zq[vX^MJNl)7�Q÷/�$�}�܃�uۃO�i�}8v�tc�hQ-��0���׾�#<�eC��Yd��q�~�d��9�:���O�Q��J��:�.����҅	c��Z20`ܿcH}���P)D9���9w�[�d�>�7�WtXy���u��W���1��]�c_��J#@SҬ|���Q�O)�LduѼ+-�����e�%�M{�N���[�8�ԇ�3w|[:�WBf��J\��5���֡T,4��Hx|&1���
�򗜉7��̛=c#��g�N�|z���P�4�{�^4�-)���>���4�cc5����Q�qΘ&���]���(y��y�]�Y��_+!z��R�hc{2)�>)���¨Q�ſOL�qϽ��\�DE/A@�E[:%�@�v:}%ڃ�\���Vhf�	���c�R�l�����E��~�Y.��/�X|�G'�\B�����l��TGFIa6=�E��o"��19)�E�m#hfRZ*	����C�����h�ia��Y�3c&�|����!܎ѷV��Zj�R��뀪7`�`�����vt0�,�� �E웰�%�On=�s�2c�Y�I�i�lG���"Tii7y��NE>�HXh1�Y�rH�}Cq� �믻ct�5Y�ѐ�yd��}b4��H�=�-^sJ�{�Ӝo��@�4��G~v�؍���!�8����7�G��7�o|�ɇ����{��
<_W`��y�^٩���V`��=j�\B��I
V+��OoƟY���56��-8~G���_w`�4K �����1V
�Z������gX������0�^�����V���U/��n�e� W)��L�Q��Jd�a���#;<�uՆ� *9�7<��䦘6ip̸���.�+���R� 8��>����$e*�Ρ<9��+"��%1��@��R͚�d\��y� {��L���ۃ�^��s��?�t�i��G֫˿�v�|�#���c�u̬~c{�ԙ��|�q�U�
n��;Xhƶ��j�������G��-��4�F���x���m��jAW�q�Ɲ�_�&�6�->�n�r^�6}
*D�q��=x��_bI�0v�UԼ޴��V��HuN��Y�126�ݛ��0�c�b��R��VT0�]na��R��2pQ��ّ�����58��d�W{+�0�h�\q����2�E�?lc��Sh�Tp ׽ �FQ���O��e^4�4������?ꎆF���,��'ıa:,�#p�R>꜓)��]�H�WBJ��u�xY�ַ�h)��#�Li?2��0�x���<1��-�B&�`�U�kj�'4-�V@Ѳ��b�0�ש-}k��rJd�.�A=��'2��y��������T\�Dz�$r���-����qG�G��w��_ N�|)S�f(��E�F.� ��N��\_�;R��}K�Qn<2L|��|�Y��	�� ^o6d]�:�RT�;��EwWw��'x��?�I<��Vd�,	h5�מ�h=Eb�_���%�W�.�҆�;Ij#'ע�%��	��d9� Z$W�F�5d��!d6��0�� �/�O�Ō�t��b!����Z�<,ݶ#��d�L��z}��9̱سk/v��/ �7�B 2ŀ��9M}��
��� ��=�V�Y+�a�U�VШXR���OmWl���|;!ј�X�c���yI,���x��܎r� IGvu��ι�?c��Mʯ��KZX�ăػu�	L�b2���>�F�e�f$Qt�q��
�[�u��b{��w,9s�ׯ���|����G.l��ħ�x1��E�I ����w�{�;]�d���r��'���^V�oن�'�Y��s«qʑ�p��>�.Ț�oX�.��g1o��u�i8�M����ӻ��5���������f��G�Ǻ�gl:0��L�5�u�^��K����@�Z�u..|�qƖ�I���˸{�^���~�� -����Q���A���v�����'8<g�G�j~_Ƹ��[�7��	��SO?7m­�M�*�$F4Hq���2`i)=u��hxnɜ(>sI��dX �����c��k�9�����w�}�Q�~�k�R�h���m'p�EѸ"��|(��B9C�ި!�JiYo"�*%,AGh�"ݡ�K~у��G �]l�& q\B.=p���k�ODL�Q�0<���;2$�gJ�8���*�J40��MItb9�H�h>o��3ZG��$:�ü6����D�R��6���HK�x=(Cc�.���f]-##�
��F��� �_�`���Qx��{0140 B��(��US�}�D�@0����Nb{u�A��KK��R�(�~�t	�2�3��}&��׬��e_w԰����c�X~�2FǱ��'��5: ���w���[o �lF~
A�)���OJ�g�=���g�G��$�M��TH;'Aa�w���G�vђ�gI4�$Ad�x�>��|L�~�L��k�R�aY�������Z9�u�2�۳�� ���x�����,7��/<��ک7�x>��!��ϋ7unϿX�i��9��
<�j|z� ��X+��b��,^87�e}&��x�;��&�8L�q0kѱ8���g�2�^�ȝvlz�1l[����s�఑J�%�I1�+��d�l 7�؅{V;*GQqw/*2�J�/���.,;l	V�ߊ�V<����`,i�8��W��7���a"xw������~l��n������A�w:�F�{.��;� ���5�˗^��t�Kট��0'ik��j���5?�Om܄D�F�n��_~��:ZT^�uw�V~��0촘�?���᳏0���jAgƸe�V�񋿍B�ԲZ���LJ �-iS�_�B�z ������HsE������Ou��o@�w�>�XL�X��
�EMē���a	0�$�ae6Թ�#N����Y�Z��r%�T�!,�L�3K)s�;��9���P�8�G&o�%�!P����O����k͹��`F�;}�p@%�$����Xd�)2���C�W��)L'2�V�PL�9~n�S�/#�\Jq"����`�i ��!f�`#X��u�fE����v]1-У_%��c�!�-J��;�c[Id��W`Z�Č���YZ����K�$ ��D�_����HؼZE�c)���{fW'��΄�j!�/`���t)��ӝ(Ot,s��DG�M��()(��Ya<d��׈R/��=��LJ�%��%�<vn&�����D+0����%)=�.�I$8��S��Q+�%h��� D���40�ǣ�Mm��|%��#�H7��Vt�s�#b��i�BX��(Y�D�ߛ�O	(�P�FP.)f�h9Z2�{�?����d�y�2Kv5ɸP��ȳ�u�"3�\K�- ���G,]����	 !x��ہ���%X6=�11�������q�p��x.S�jj��X�y�*��̡��Q5l<��F<�f76�@��;n����N[����l ���X&w�\�]z�y���g�>�A�~	+Ě�>�}�7B5�Ҙ-�Ô�0�����隉�݉�=�+w�Q�]pD��`;��"68I=��8$5���JC!O@�(���!_��q�Q�Ek��|JtĐ��%xwd����՗/�
{'*2h�z�a����ǜ�ܽ-�<R��R,��k����9���E�I'1��6���.���݂U�V"�6��o,k�i��Z2��xtC���/�����_������-e��;c���c_�:�f���= ��@�TL'G'(�3,aϟ�5�L�jQ�6���k��E֓�H�`��� h4E��Y� !�vPSO�D{�	xy�K�WQ�A)
��	�a$2�(:JW�[���@�����Pt*���%�-v/�ё��i�Ӱ��[
��h�1w����O���T:�j�=_��!���QI�)�&�6��tbTS�	I,G�8~�v�><DK|
���{I���6i�4�x����%lz�dG%]���x�1آ�9���OI�A�e;{�^-q���?�'�R!��Av��׈�ji�%�r.����FF��4�d�A��㥂�5,�� �͟�G��J��J�q)M���Cخ�k�77�8��M1��*��X�]@�Ϥ���kď�`��r�~H����p�LE�1���F��t�S�	��U��P�?�|���"�Ŗ�yq����Nrc�A�?�Ȧ�3"��!�]�[-��K��������e"���|^$�>���5��$�x-/���_%��b�7IDr�k��/a���������
tg�8r��@��=���`zw���X2�B<(L���w��o^�C>�߼�S��Ϸ��TE�?�L4�$Y��<��G�h�)i�uZ�&p��,N�߁Dy��6�F&�(�a�a'��Wz "�WEGw��}��_��e ��cr� �.��冔��t?�FY��&}4��ѳ�`�.��v\�0ؒ́4Ԑ0B�!��"�锆b�`ao{�+��_��8��B �tSaiW��<ZT�fG͘nl(+��K��Sw��
q����b7�������'v��ϙ'���O9��vaQ�3Q��zh�����}۱����O?���2�.����Ү�/|�#8��~�-ݪ>�寡n���R�Z�]��e�r4�\��F=�
��h�}���})�ʟ�Q}���@�a�]h�a�P�O �IC�=����iL��`���s(��Sҡ���;�����\�'4Cb���t���8B(Qb"d��8ߓr3�o6�L%�	��z��D 1�Gl	��L22�BJ���X�j�,�S�.d��kْ0�QPv�Joh�����m35R��i:>zp�}�P��B=��eo�s��x�MF��E48�X� �(}L��P"Z	���O3��\��kCiP�^����Zg�6���t���?4��ufi�@V�i�M��[?#4N3��Im�.��I�T���i��t�uuc�c��a�i5��"�} ����Q��7|&Gq1�{��W;s�q(Y7��ᚾʯ�㱷|�=�	�jy����� 7k.R]��_(��/z�{�����a��x#2��V��$j�j�K����b׫�y���{4Ҭ=j�y&�A(&�)[I]��o�P��m��a�:	�f'�M	#B�N K��������&� ��eL!Do��/���1t`	��@.�����Xܗ��,���r�����6?u�ϑ�zx�#b�0�+�y�U�5d�k1��8Y�w�X��cU�R9�)G�W1'g��%�8k�4$ʻ1�s5�VI�V8��Է\tȟ���լ��ٙ~}�ފ��.�M���vt�Md�W`���Ht����*JH�@�@%�В���MN�@2�X*+��^q�_Cڎ� Q��f��5�R��6��Ⱥ
lf�5m A�����#����;�c�xY-���oΫ/]~�|P�<~9>��^�ER��G6��o^����� �2�x�_�O�{������Ld~.a��Gգ=��_�كk���R������m��a��{�9��y��&ղ�.cŶ���O	;��@"�j3�˸T�F��t�+������7���#i��w��]]�ퟠ޲��C)���\j�I�|��?`��SG�^��t�fi��J���ܥf�O��Q��2aK��tDR.I�5�h�3hVpR��4���ʡX���=�%�����L�H�(	��R[�����G�Z�kr*&�Q!2ɔ &2��xR�+�����`�_o �����&Q+V��Ѻ��.�*��/��nM��_�N[�P���H�x>���'�jq~�
�xb�S2}#�+��Z&D6P�ݔ �	��y���7Q(NJg���$R�Ĝ8�cy �E<�IQ�M�x����u���H��1�+�H�S�c�ܹ�鍿��K�[���ƐKe�j�j�������{Ou
���N7����a�`#���Q��t*F�>,�88�]�	�Y-�#N������d@���#{�X��0�hD���Ar��P�'���=te���	��q��7(��@y����TI	y������I
����^��_���H�7�ݓ�K�Y�P�|NG,L�"�������<7:h���@�I:��y��\����=�X4w>�mَ� ��L�|�+�P�u�i���ύwƩ��Z��
L=<��5�z��زs�������lX��ܿr+��`v��ĕz=��S����Ӑ��B�߅���j֤�:�5/}��n=T��*���G"a��?�
c�1��%CY���A��!�{t%v��������&����Cy��:��s��YhC�����h5�FG/����{e�[���\;ag���&�$u2!u���i���ԛHY��!~�˫�Ϟ�G�W՗��6�=T�u���p��o2��Z�rcx���%�D�I#f'�6K�x��G���i��V���}ƶѺ:0�����9<��t˚_sۃ�+���3��g?�!��_�[�C�����=+����E=л��-xN�tRz@l��Y9O��{��e�lZF^�k?�����o@+�=?8�� ���U��e���6 �A��7Z%���.m蚁ş@o�d=ƍ���ve`���`�@��U��0��`&'%�,�8rǸ��KظB~T�Ō�RLW�V���A���D2	ۈ�R*��>�`9!�u��dR�B����I�8���'Q�w��O#Y9�s�c:VaC�Gho�f;Q*z"z�\[o~���s[dX:e���
Hq�VMtu���Q݇riq'�7�}-���W�L�/�BV�q���RR�$�:���^�j{v햁�8^@��K���ٰY��+;�v2�P@Ϭ~��g ���{WI�<�J�\)��09���G�+��J,�;`�tσ��3�Ӈ'�Z�5�6`ێ=س� &&�\@`d;AS�t��&�	tt��q;1Q(à'����hNͶ	��F&��L%K⻐2����R=�=:*���������/v�wta�'"1}{���+v,.�S}�J���m_��ȼ/��/�ŠY^�{Jٕ#r,mNoS�t�=��l��lK�! i+��h˦e]"	$�A?M[�(������x/~(ɴ�b��p3�?7�׋y3gc��-(�j��Sq���Œ�� ��_x�!��~��7�^wj�+0��<���1<gV`�]j,_s��L�~lۼkv��N1`��:�2�]Ѝ3�@����L���Ĉ�ut���Fv�!{�
c��`�|�# �X[�8�4[��^���ˠfub���002ZB+diW���N=�vNg�.�F���?�#MC<<��N\�?�Ф��nB̿����q4kU�L�i�b�w��G�a՘R�����W116�7�u���o����+�qG	���/c�	t��m��GЗn�����}��c������_��/��׼�_a�3X�`!����pD�3�-~��]�s���ހ��i�%����mL��8�����;nl����icˁ���g/�w�+��۞r]$��iC{�"��)��,q�c�����$�0�ʠ�֨��Yv�L?
"�Q׆l����(��z�k�p^[��{�2����~-�"��9��}Y�KcX�n%P�Y��^k�Zv����L.��R�c���Utvu�#�E�\/N*��`�B�ܷ#�I�vQ��6C�ar� `6f�E�(��(��`�����L����__�Ɔ��7�t���:I�� �I��j��+���8��	�ܱ6=d'�󃃨�-����h6�DWW�� �s�^gٜ�Ï>�R~R����~�;��B'�vf�Y�?�|+�|	}���.�?����/C�0�/|�Bĭ���0(q7�ys����01���<ox��	�    IDAT���O���uc��]Ŵ���v�&�Y�N��f����v>0<��c�� ��+���XE�_*�`*쌷�E�L���6|tի%�#��&l�-@O<�{n�O���ӝ�jM ��oy� ��ɼ�тjS=�U�7uW<!A��n��&u�|J|D��=2���4my�\���c�pA$s�������1��"D4�k������2��%�鐍�26�0F �@f�c���ؼq3*�b*DW����x@lo/9�C���9�8u S+p�V`��9D;����+@�x�(�H!4p�cO��-#X�sL�'�H�R_\���rx��s���@�]E:�@ylAÃ�����8���C�����c������ګ��)��mje����+Vc�h*5�0��0�=�,����J)w#C�0Z�u��톕J���a3{pͷ��S���tU�\x)�X�-+7�%)�-�'�D��ёH�����IX�<������#���/���=	�V���>������R��2��} ��>-6�@u��_��G��'f�-}���52����?�cK���;��H$s8��#p�O/�_��_����_�Ju��Ch���Zr��a�^z�r���ow����{��E���[�5� .�Ÿ��}9̝щL��%�Q�?<�r%�j���8�\\�����z���2�R6R,��N�xnb�xy(>�ݻ����P�]�O?�َ���0�>�,��3�:��(V<r/ܸ���8N�92 1�]� ۷l����q��#1�?��]�3a��	tv��&�:8�ēЕ�	cdWoڀG�x{�GQ-T�?o)����XQXʄd�[X�(�Jv�9�Z�6p1щ�wؙ ��G-ݑ�z,l&V�Еˠ��Ų�pb!�ŲH���4(�DU�Vt˃	�)q-�.�b(���y������c��A�����$[~^��S��_�
[7oC:�Ĭiӱ�E8春�̺?�G�i`Z�x}l%n���5�Bs���	'/R�j���dM�=d��vt"���(�R)����>k6nބ�[vb��Q�S=��]80Z�*�:mLzkb��!����/.&x2ec����u��	���^]�u��~������@+�����X��o¦�����Ѭi��x�#��O�&�^L
�x������� �_ˎ	�؋���,��fC����>'�џFV�m�:��ߗ�1�Hf�:L���ْ�,�E���P����������Ad����M[��! y��_/ đ�)�?�;��Q?V��Fυ��:�������[D�ō;���x`�F�������BC�oj�����僘�*"YB�FFȖ]�zۻ��#9��<kű�*�cE��=���`#�R1���q�J���D�F��4�4m���)���g1�2� ���&�d�\ӛ�*��݃뮹Gfc�xM5��x�U���UH��$�1^*ˮ"� ��$z;�ว*��<n����aca�clk)��K��}O��p�Y��;��cW���d�a�>���ᱭ��=k*���u�F�y��W/�K��Țn�P���]��jN��7~l��3_�:v�����`~Tt����>�e����A״����ժ�>����[߇������>�?]���]u�o�O��ې9S�����W����?����/ ��?�x6m�,��Ԩsw�#�ìY���π��A�+���btb\^����w܅�bf��ٯz���o����ibrnzN;�D������ǁ�1�L�P��O�X����xū���m;��Ï���G"ב�5�� 5��z��?��(������-�gvv��U�B B�DoL1�6�0`l۱���IHp�����c;�O\ƈ^�꽭���vW�����{�ν�y���j%���.3�]vfn�n{��}
�u�`��/�}��6�}���_\�
^x�U���F���ֶH�l���fq�J�h���h�y6����%��"��R�,F+Ԏ ��(d	��%2���hoA[s.Y}N[8�L�KCEE%v���Y���`bb��.����oԽ��X�����`6�"a?���JTG+�u�V�<���$��ZZg`���x��0:4�|V�T�P
0؜7�W_~1Ba?N;�"�W׽`�{�G����܂��ZNonm��� �{�38��|�����hjl����:�?���y��v�C��!Ȟ�~:�HgI��r���E���B0ݼ�h4��=G����0�I�|^��_�|���>t[�o���9�A��{��c�P'�j�/�,��D�+�$q�s�o'�%�F�XA\K��hFVǥ\��6�kE/v#+^���#�e�8�N)�,ptS�E��ݹHN�*6d7�_`�HH8����i���*K�ɂ�@���zt�B<��v�Oş��,h�S���N�r_��>�ʟ/����/�?ģV���g#�m�A;���v���l9ԃ_���i i��Mnr� I@��1҈�m̬V�
!T�W�DХ�--��#Q,X�-�C���6v >�i�T��1�}�l���#�����`2[D�P0�U�,z�7)a��b��A��QP�,5	�if�mFH��Uxd��~|�<�z�;')�ٓ��g֣g0΅Qޒ9Y��%kU�d��J`��6���5�皳��i[���a3������]3W���/Ə��/D'#]�_�э�~�KH���E�09��dw����ǻ�;��r\���-�ak7���/Ea����_�ukDpر����V��g�l?����� SYhF�Īo�s|~������sŶM�m���}���c�BvWp1��e�IE��r	��m�i�1����}#����v"�d[U*�|N_��-��u�m�,b��x��g��� �ǎ@�z���������y���2H	}��ֈ�/\�9��1�ׅ�C�Y��J���>�ÐT*�+��܂ys�0HH��<����T�{/N�3�������;���c��8�9��UX�a7
���!:$,'j�Z�؞������f�B@NM4�M��A�4� T�Zd�k3հ�6��+���%�q��bF�	�I�姿xʦu�����D,G2����0zzz���u�y�jY�d:Z[���10pC#�ط� S������y&l�L�K�B��Aȫ����J�X567�c4�ƾ}�X�h�]s&�H�Rhnk���T<����� �Α� t�D}}=n��&�Z.���>���n�ft��|��yd�D7"J�9U�+UUDX��3�_\�[��d�XȖWu��rU��)��t�\�5$t�Н35\"ٝ&M2PD%��JA����kq��ZQ��E���"������mW/� ��%�Ĳ��% ��i��['�a��8dה���J*s����V8�ml�%��	l ionFwg7������_�]�^�%-��4.9�D��x����9e �y��{�#�e�~;_���M� ��[��Mqd$�����r��<���:�<s��!r��Tr�	��	��Ub�5�+��֮�t�Ƕ�,!Vb�6�����P�wcbl�g���J�����=5؈����/vw#��>`�[�2�������Y�p��d���Y�o!�IcA4(�z��޸������$(� �y��ǂW�ĸ�pŅ���o������r������/|��W���]q�\���wK=ɴ�
H?|u���Y%��䁩�̺�����@vl������[��I��K���Q���Fzn{���=��Fm��~�_pz{���>�a������mH%s����V�7D��R��o�3���3�`�I[�X�e7?`���n�a�P�(5��Kל�s��ĕ���9�5oy̟���u	�n��K��9��c�.*���]�h��w_�M������_����Q�Ԉ��Z}o޴�����H�Օ8s�R��6�y�3����Ex<^���#��9�����ȑ#���L�����O��k����L%|��g흻���?�j��p�����_��T��\RW�.�(K�ƈ ���!zUsgq�(2R�1���B^R9a�P�XH�/�4vJ{$�s�b\u�J|�k�0�?��6Qt&	�9�x"����������Z���a���L���(�o��t�H7R�:;">>��KF]M-�)HО�f���l  #��[��!��|�F
d-��Y�p�wIC�{��a�~�����}6�k'�)9փ�1Ț#�cL!�袋p�U��~��|�~n�zlغ��ꯄ��H'Eu>zpkB�E{r�r�!���(�*�]��Z��0�)G(�R����8"˅�srrs�S��\��;QB(�hA+$x��N�u:@�~R8�tw*�\��k�A���^� =N3C����%����ʓ��^��:k��B��;����cA,�TF0w�L>܉�x�)X��y4������2 )�x�#�[+�����W�ߧ�s�{
�dM�ˋ-����82����Md��Hf���y��pI3
;Q��Q���A8�n�0c��X��<h�o=������^[�-x5wlB�^���Ue�SI��$o=�xmg'R��Z��T���G��r�&����T(�t#�
�8�#Td%�\�G�_��<i�x��$��y�J�}����a��KI̾����o�w�v-fQ���1���aQ�_�ү6�?�=��v�Z}�����n��v�"�=4f�o���	��J�M-��65��GA26��n�	���}oz{�kľ��wr����s���~	s���i�}l,g�W{yGl����*�p�	`�90f�Ⱦ�*ğ{�����?�i��� o�P<^��Q���W�/�e����u��m�Ν��0�9��An�U����-ܰa#kZ�Z�+GZ���ÈO&���`�.��9T �bq�^ �uKS#�k"<��s\@��A�P&��rJ�3g.��LҼh*�����d�?��z��>��}��/���t��k��6.��:�y�G���wAR#���+���d�OC�2�'�ߏ�g�OEY��m�]6�&T�}q:���Qڱ�ٙ�����ӓ����0�V�;n��W�a�֭[o��Z�\�Ǐ�Ǐ���&,^�g�<��enM��Ӗ�%��v�c�#X��K(d2�*<��p��ԥ��c[Wr�b�U��t�P࣋-�Sd�����\Xv�yX~�ұ��v��#pPa&����(�G�~�&�[���a����p�"޾��}ز}�z������)��r�J�H�b8T�:I�
�<> NL�J�BKdN��A��%ʑӍ`���A�TN
g�PB��Y�Vq&=�;/�!^��R�@ps�s�"�H��nu����O��Z���WhSN�zK�{C:��[���Y��~4�R�.�2:�$(���HfΘ��|xhL�܈e���8�8�����>^�ly��G�@���~y��0@R�b��l���֮A<��~��#o)��
4���բ��Wʢ�m�KN�<yUj
�b
%h�|H$3�ֵ����?{��\&�m��^.��+�o�6�tD6>��Oc�~^7`�=g��H�}	����.�1���;0��!�&�*6�T[(�D�r�
h� gM�,�b��{&���\��p&B��L6_�}�Ǳk�.vd�V�rq6>>��χ��碾.�b�9U��h�{���_?k_~��
��a��ҕ�׿���!D����c�e��ǋ\&#6�d��3���9�Յp��w�7]25����f�J:��n�����͙����w4�G���3������!�S��<���;ڈ�)����c�V�������w-�^���ۻ��k���={&S�����Gv�_�;��"k*	����1u$��#�IC/�9AB�T�ܴ(D�EUU%\2%�������A�ZH�|�M���2�HU�g���v�ލ��q����k֬������?�?�����/��'\�3ϻ�������l^Bj2ů�̧3D¨jnAEu򖍱؄���SٲPW[���:�L޿{�7�5�����T�<8c^���-���7r�w��m��F,c����(;Q$�swk��Y8c�2ؖ��i>����}�t�X��{�ؾA������aM^�������D!��B	�x�m{��V�1ν���c��?<������9�p"����痘7!�Z�б��t�H��d:�D:��6lBEM���L^�a����=����n��0/Q�Tց�BD(�(�E��� ��7�0)�K��w;�T��p��Tnǩ.V%Az�z� ��2�/�wMD0�tM�^���2���q��'��:�\"��$N�d%L�O�O����(��X_���H�-Boo/�zYv�p��o��Q�������R~��G�<Sf��(�@yh�w�I|J��I֞Z ;�����=�����
���f�L�Wv�������q`b ~d�Z�D�\ք���r�hl�	*!����W6�c��/�.�d��$�8�oF{��U$�6�S*@�'3�<>���V���u���36�&�guؖ*�4p��6!!g(W���ղ�\���N��.�{濱,$*���Y�
���0f�$�3��焽�ቬM�ZD�!P��1(=������/l؂44��R F.�����!�:��e�ŝ���~�-n��,�ꑧ4f���� ��ah��+V�����Cұ���^���G��1��'O \Q�db�; 7_��b���̧�N�rx蟾�-�����ti��f�,�)x	*p�g��+�ǚUoo��i�F��4F$<�sAT�� z��O��_���P�A�d�"H�^E���h%�:�oT� $�/����&��O�3p��>�:��~�Xq��c�n{xl�úu�~ë���E�"�ݙ��<�,a�B��{��?�����ӿ~�h#��z�Ӱ%@B~�fK�����T°��	�+�
YD%rA�dk��4(�ۋ׬�sk�b�X�Hæ|MCȫ@�2��5����ca{�^C_�j��Do�qv�"�)Ҁ�ho�����T߀5�ϓz��أ�#(��!a<@t�ʀ�<��;:�ѩn���<м�U=�e)0�"q<u��eX64-�D���ހ��� m[���0`�x��{����!���O@��8w���f��~��$��7�6�{ϼ��W���I���⮆-�!��A��+Fz�fp6����]�)���5xcG��`8�D�"�Bb��) �O)_p�k�t@�
�L-��;��2��O '���F�4�S"B(Eb	�0+��A�2kN�^' H�-=G�e�"��i��Cw���UB����5�~�{�or�)�<j#P�x�Ԏxy�v��G�'�*�vi�Aîc����;07Q����M��f�=̍,���5>�Z܀-%9�>�ư��f�Et�DMC=Zf�Fc�, ���@���8=����G�
Ǥ�"��8b��8އ��#��Evl!nz���e7��9��g8�d�����W�Xޅ��,�&�\dU�B��`0[�qd ����&�[���U- ��{n�g.[��s�qzP���flM�af���@���w{�U/e���p
?��/����H6������Д �B���sW`��%��E�}�9�ܱ���r*L
�"y�
VI�nd��ͬ�* �u��=���̋��˧_�D���=�f��ˏ����k��D�n{���Q���F�'6i�UF�����V[�{�ŷ�^�a��*d�6,�_PI� L�*���<7_�_�������}��a�F�������x�|��}�o>�T*�	��ãhjja5�z�\���s����4O c"6���z.Ҩ#@��R��Xp��'>�ŋs�%�ɣ��[6o��[��W�P�5UU�MK�,A{�����6m�Io�����v���-F<�)��}p�eL�r�����KgP$!4�6<��,�TWF,e�	�S�6!��4D}.�ǻqř�����e���H7�v�ޥ���g����G    IDAT[[��p�B474���3�gH7�j��� ��B���Z_���N���'ǝ�m�� Ե�{���b��n
uY�lA�)�x�mw���op Uu5,�'�3'�K"��G?�1��4�:k%4�;v�f�3r�Z���{m=��-Fg�6����.��}�\��"�Qd�[z9t�i�$N,':��=��!�S���rE���ą|I^�,�37�[�Naqh�ӶJ7^�|�}G0.��(l��a�4'GdJG"���W�c��Y�W���'���Lt�?8� �s�{"A�Ty�uc������YF�- ��uS��ß�wv��*��x�#P�x�������9�{����,]*R��}�cx��m�P��E�<#OE��e�����X�^��D�*�8��a�5aM�O�9܍Ҙ�g Z�������z>υ �<T����L�}��?9:���8�l��9�S�(SA�p|,������+((Q�R��x����2鼠l�U��-��E%!�����~^.�:�hR�c밍4͛����U��\EC�!�*�h��8���v�$=ם�����c�!�$��BxB���u��;��$�b��d�;�7�<�l<)�n��^4��в�r>��
{��'| g,]�o��������% �(�\�<.��b��g�Êia�G˦�g����ڇ�iR�;����[��nh�0��#���^	�a�*�C�
���s����d�ҩW�ƍ잾�H&�;w.�~/�z�	ѩ�����f��:67�x.��R������y���䧝v:�9w�O>���n��F�Z=�������J$Z�����3g�d�b&���رc8�롢��X���V��zc���K��'�mÞ�QX�&s�ҹ$(XENLGބb�`���^�4��P�Av�"��/�G���TfE������9MU�?�p��>�ֿ��㢖� v�����$8_�`fϘ�sV�%����C�fX��V��}��R~�������{�
]�*B��zӜP>:��S��D���K�p��7�.��|���8����76��6�G�������Nl�}��1�7oV�Z���wc�i�10��~���������h��P�.f�@�%D��g`�У8-���igi	�8���c� �7 �R��)'�I݉��Lm��V� ����: % �ˡ�� %z�`�|Hp�
<.ꫫ��ڂ���ct�,�]@H�N ĕ�(k@�8ˀ�^��F�@~G]^��� YDe��5qx$��<���tSf B�~�fI�*�h��c~k5�@TI!h" M"$����*��,�䅤�!|���g����� ь-�d�I�sC�!�N�ؑn.�2�44E��x����mT/vu�p����C��"c��G ���G*C: �n
 � qħ�`����oޤ,*%U���a��m!a��X�p.Ys�*B<[��x�4��)a���c?�RAR`�1�P(��N��,^��s��*�AĆG�����b.�.Hł [�Gi�ds\�L����[Z�008C/�*����Ӌ��1{V+V�X�e�g��)p{d��&n/k#L�`:���~f�g���x���8p�(y8"��	�\��Z:>}�p��_{o}�W�=ǘjE]y^����C���{�V�Z	E���{;��[� eΜY�1c����~�~��_q��}�~�������W������ z�!l߾�y��u�TVr���܇��Z�I���T��q�f֦��`&*֜ys���t�R̙��\�����6�Bo�D�R���X&�+z!d��/ŒQL��%KN$�S��Q, ���Ph�Pe3�#���]ȡ�҇W���[����������2%lV���C̛7sg�F�*�l6�t&U�O����ʶ�m��̔���?i'G�a�@�!�:KD����#�����*�n�(�	@�|x�o8���X���0�~�����s����/�{��XEַBuc0s���K.�Ͽ�j[�Q�Cx�ɗ���8���ދ@H�4P �'���Y� \�JRD�䋽�a8!�~�v�t�N����:"���_s{/��S��{"2BD���@ћ��iUԍ/הf��Sһ8����Ҁ8/�" ¸Ķ�)
T�F]U3��p��!����P�����p��zX�\���_{��a<��[Y����/�������{<$`&
9�.�LG&��?/l���r��0�#�����Ȗ��Q,�Հjwi ^sU�<�,jC^�(�+���Ԥ��&BE	���&�]ۄ��r~���BM~K�*\�K�Dp<G���k;��"�V4B�Vch��X����qL$��$��A���N]�`��憤(�!��,d%��T4�&4
��TVV 6:�%�#���-��ɗ_A2�����y�B���S��4 noFVP;$��z\�h{
:R}��A֗�O!�U.X��|���!jU
n���/��#*B�ۋP��h����\��(*�*��o��%Z;JO碘�nS����zB�&��(
�-ܦ\*^�ku������G~���K/�`���h][������aA�m��Ɲ	��3Vcc���҆.X�ٳ���o~k�>�����ߍ믿/��<��0u��G�s�,�n����$.�7�V��(>������p�
��~��Wx�n��1k<>/*+��|�
̚y�~iog��i�A���-��3���N�ڔ��H�Nי"&l(�"��D>��A��!��WD0�J��&��H.x(���rYh��?��fDNU>���Ͼ`'I�Oִ��T6��LA��X�hf�π���d�q��]�e#�I`��Y��£_�*�����! յ�$OڦᒌҶt�������yC�6���{1c�j>��jO��uG�h5&�x���r�il"�P8�� {���܃�u���o=b'r:
Z�{}��r�m
��!�4_�e��Z�V�v�MJ.X��D�qeLO"����O�+�N`27� ��]��$U�p��=��\�� @���(txK�S��� @@4���@E� C��#�wܱXF�";�L$�h���t��%���ى�G��q���&��z\�t&��.=�D�{�8/o����F���}(o^y~k#�n�6ۥz� ϚE��`��!<���'a�l�+f��v����B%Ѻ�gMHuHC{�Kg�'�SP�1��dD<2��&�y�T��j�S�|���
u�R1E!��n\����c"m��hY��S	hQ@�`"mb<^@��[3����͔��}Ȱ0s9x�௨`ڕ		)��U4��DϗX�LN:�$�Ҕ%@�hD��ɖ)<�I�
Z�I�>�T����"�T!���ؙ�^
D4-�ԭ)g^ 1�*B�(I���qh$��]�a��E�V �x)���e�
�"$�#�� ��w���m�Ƅf�-��M�^`L��Ρ�I�o�E��u?�����_c�����[7o�l����hB�͘=k
�#�@ ��N_��q�F.��N���R����"7�J�?���p���=(;v���g��5 ���/������w��!�A/��|������`5Q��^/^{u=zzz
W0@���ky��9���$rF��q��Q~Ȏ�{!*��phpI:e,C�,,�bQWe��%�t�����Ź�)@r�g������nz�bE���ɠ�M`?����|�cw��3�h�pp�M����s|�������GI�D![q�|�yC:�d �ukH:��GC1��?�/��8lvT��c)(AT܊�]B��9�@���P�|�����y0�ĞH�161ʠ�,��8н��?���8k��Ҽ�`�۹���E�{h���'�Fnl�م����j`�.�+&0I+���iL����!�q���I���]��7S�����Ś�7ÁӺ��_���ŴŖ4 tmN�[O[>g�L��)�W�Q�����t:� $�ߣ����i�u�����M�O�Rl��l��P���X����-/�Oq� �O���-G`��6T���E�rvƋ�{�5���|�ɧ��.��BOvv�r�db��'J;*��i�Q��u��<�$j�*��
�
	'l2�e�5 �ep��ޢDz2Q��y�-	�M	���T���4��L�E�R�(
e��g
�H`2�C��0�˟�[�&�l!�m�'c\ ���ŅX*��٭1H�P�Mt��\DPBE��㨐g���%� ��v�6gy0݋�KI��Ǎ�Hz>�b.�9��PuFbB��P�@���'KT
R��@�&
���]ԩ"��<� G�L� YbV���,@)m[�*�Wu��%��`�IN!'\wL[�GSA����~#�G��o�z��-��:�^���s`$��������MNk9��Tᓟ�$�h��g�k��#�`2���-[p�� ��ك��f�w�}��+�����w�6��m-x衿���{���@��R�M�zi7>���ҋ�����n ���u/��]{v��0Ee�9�Q�؀�����%�WF�������N�u�o;���)z`Inh\�R���:h��z���J��� �x4�s�j�Ϝ�g��lyr=3->l�\��y�U|��+q�%�b�̆�q�9�kS��P�aN'{b�b�������z�j�<�,�O�B�.dAg[��h�i­J����^��/���X{En]$B�N� �䘥1��M�F0��T�^��W�;DFM�m�?bW.��9I�TV4��'?A�`"TFMmI�"���҈O�c�=�3{�}����ы�X����ӥ(�E�$���	���	��:%�oٛS�J7�_@ފ��v �:2��1kC��X�r�>_
t�8}���t�� ����k
���Hq�{ַ��d��P�9 t}%�)�xS��;ލ�fׂ �U�U����Dy���/�w8p��q��k��ضL�_�n���-}xiO/���(9ə��T��G>%��C�f��\0��f�U�6��>�FH�!g��2+@}�j1���.���z���DsA�.���H�i��D�`2L�G�XOPU�H��<�'���62��H�X$�/��.�-R��f ܕaԵ�0�%k�$i�����1�c�mF&v$�E!.yѡ2X�e@��M��'�-�~���
�Pв��e�`䒰&ӘRm$�u)J��p����.�:"�]�D��H9�(p�(��1�`pG?�uA}%U3����zDj��.�xB�����*�-nTT�hR�B���o���".^pr����e��v��s��O�˂o��lt�%-�
�|5����^�.����KX�n��b�ޅ^�[n������?��{�?��҄O����r��>l۶���a��L��5k|�A4440��b�hK�_Y� 'RQ�"��s��D8�P���Aoo���d6��t��`�#(��.Cq{�H�|�*�P!�������s�(��BcC=�k�q�E�� W:wٚ��ԡQ�_1�s���މ+/<Q �ر�&����� ��HD�q�8t��+#a�s�9Xs��L�J'�M�qG�����y=��mP����|V.�p��|ޑ�i��"�?Q�XP����%m�܅��#w��	�L�Nm�W����|�;��Nu���9���(�������=Cc��ه�7�E�@^>W���W�*(�ԏ፥���
�RJx�UwZ\�oxC?�#rB�QZ�TG�q�*u0���|�:/t��=�Q��2ߜa� '��t�u������T�Զp�o2Sv����t ���� ��'�����o`����+��k����)�<��@��)���6�v�I�LE�)�0/^�q�m�b��%sF �hv�(hFTl�(]�t���P�L��.��U�!�Au� �c��4��C@�����
��L��X��'��jJ��Li�b �/����BQ����F�`�i$��Y������E3����g�mȡ ��QX��4�-Y�)��s2Q���(D7!�.-�d��Ќ�C�hS���ó��q`� ����W(�]�#��d��̩D6����l�F�g��E�$$AE1S:��.��2խm� �$ۄeP�6$�X���Iu�B�ǆ�+%�₻�
`Ɏ?��Y&�����B�gri8e�@ͧ񷟸�_��3��:��\>�ݏ��,>'�+*>I@��5�:w�y'�uD�>�l|����Ɔ�P� �	Ѭ�����^|�yTWG�8���<� �;���O]���'\X��}�ß�ٟqL��Ȣ����_��͛�'�[�Ѫ:x�~-w�X>��Z>�Ś!�ri�(�Y@�l��"{e�A�K!�fr�쭫�!�L�jlnb]Hj2��Hz&���!x�\����1�B�DE?��nł�C�k���I�y��SϰW_}ͦQ�HB�zI��uvu����īV��]��AD#Ȥ����H'x��G�2��ڵ��Ydqv�
V�yytm�2�<S�;�C�A�i�%�壟��'3��&���\�5822�����f3�0���444����+�O�d�G�[
;����9\��E �&�)C�z�x a��7����ϜRr��S���c:��
'��:���w:�k�W���@��� ��� )}��Ab�b�`
XL�Lw��{�I�2��RJC���)X��hind�d"E�Pl�}�X1���$.=�rU� �#�G�|�Á+�s��?l�r������-��̖�@H2���L{ ��Ne�,��fy2�2�GUPC{} ����dġb��ښ���I�}�UA�b�'UɊ�D&ϓ�&�L�]�|�z�m�'��%r����J$���D��P炉[ 2L�&G\���V���VeL&���R�m���P�M�<�(��T� -�pSĠ\E��v�E'��e����T��\�vEqlA�B�Dzb��%��@���ma%*�T 8c���^B�m�Է`2�E�ȡX�@��P�d'�HB��ҫd/J˦��D��`2';��dg���R�D,�u�|b�K�8�Z}��r�p�AH_πM�cdl��F@�B�&A]�{;�d
˗/�g?�Y�q��?>Ȁ�(E�������M|��g�V]}����|�K_�1�GsS+�|�O��^������[o����a@% L3��ަ-�Q(�����=w!*��H��`N�p�������a`l�3�w0I������>?�Q���5B��(>k4\E�a��T7w��L�,Ґ���Eד�vs��K�$=������g��.�z�����c1�#�	��|��E_4�D�J�c���4TVT0���G���K�x�gY���O��)	�������2eRS��fq��(X�'��N�M�;�ںe g�`�
�
���8����	8�VW����d��|CQlܲ�����j���QH�!W5�H�i�n���B�x4\t�pވ#s��' ��~�����K����YⰔ(O�N B��	��i�� Ƞ���t�
�S���; bJA�����I�4NI'� U�e�{�]dS	 ��5���F"���J�z��[���z�|W�sF���u'I������/��Q�i#��`�M�>�:e�ˍWvu����4P��ߠ��	#�D���"���"��g%�Z<�O��U�W5P]�!�;*<*}�~���l���<�ؓ���ķW=~�|���R�l�	v���L.-[�d��'��H���#t�\��������Y�@"��J�u+����`����
�+*���`A�-��X3l6S�(`ML˶�"u��y!3����T�HFzl�g�鈄Ɣ�My�@��F����-A��T���r�סu�LR�c8�A&��ۣ��OBʧP�ǁ|Qϸ��{D�c������f�    IDATsӜ�h{�����������K��	hR!S�#$�����O����t:Ʌ�}�y�)�cƌ,B6
y �"s��Q���Tr������G��k��e�X4��+�`߾}l�+�;�L	���O�(��m��FmM=�-=k׮ePC ��#uv�˳�����b 
����x���M�������?؁�6n�'�h<���Ł��36<�(G���e�P�^0tq��5�����"0�i���	QLS*o2}J����߭��i6|v�ݧp�U�4�]�G�>$�iL&��q�◨l�(�d��hii��YsC�gA��\��6�{�Fز�� �h��'��4D�(PD����0J��P�]=���CAUC��'@�`����kdxLM����?���:�#�9`RF:�E���a�Vtt�B��ml*�1:8�@G7��)�p�֖�b�- �U��3 B�'qݝ�S��?׉�	����L�S�T��� �P�IZg94�3�^I7F���8@��C�G9 �Hl"	�WESu��UhKP��:�L�*�x�#P �t�����ꀤ��`����ac�1<����s�nl,�N��u�#^$�� ��U%��gxV�[v!A���P >���l`�-/��,�ܥ}�KE:k��m�S�`"�g�O�@�����(��,����1q�e��0u��Atf��
�Ar�0�Zt���m�'�N��.���+�^�G&�����PT7,���c��U�*�\���[Pb�C!ꚙK�� �|^h4�I�\�$�&%ϱ6��hPl�<�����5QT���x9��11���� �,<RAم��Ð�W�Y>�=H�;U���T�$�C�ĥq׆�k��VIDOyd�,fN=� ,�(X<�y�{qÕ+��G���|>��u��	��`=Q��/?��H2g�A�S���o|��PtNQ�5W��>�,v�܉ Y��2b��x��'�SB�fr�"��o}�hjj��Si׮��������݈u���'�>��}�k����Ýl�,��9����?��[�V1��5s�5����S`aב^l۹Y�D"���瞇��!;���W��aMw��P�X�s�-�a$Z!9v���!�mQG��-E�MTɂO��G��=��{�9�v��ۦ�g*�D,�����OU4�e˖����u2CSC=T� ��Xl!��\���s8~���Nd���Ú�C&M
Ӓ�Z�WA���:ՋT�Bư�܃HM=z���g9�qbr��i�o�׿�M̜=��#PI���Ӈeg�����/�����
w 
�S�<�-u��pҼ���@���Q  _�aq�/��KPEK@����kzq_�6~�M�MH	9����|�K���&�'�-��T��UJ�u%�`���j|�p�Ka�@���kyڸ����#�t�����ڊ]�vadx�����x�MWbfD�jL�Ue
֯?Gʟ(����@��ό�L��{�Y�p��m��p?�?���#iX���d/*:4�F�BB�2%�Ѓ�:I*r�ETz_%�uL�!ʦ�`7T�u$�rH�4E��I<�M6��`��b�f�-. u��ă�EA��a�2��
k6H�~����A�<*��J몐��r��*��i+HXmu�^��>J��*	��ǇȲ�6
��s��G,�E2������<���7��e�,� ���
d��M��߭�0sD�NY ۰�� �!�4w�0�:��j��j�+�C�X�d*�b�:���2)���d'����O��Xn|�ؐ50��(ZTTRm���l�+�T*,��8|��U�ѲY�MԶB�9��f��q+�s����-n&������a���a��3�1� �(�$��O<�w#h;ɽ��|�uԭ�z���x�3`hk�'���36�1�����Ϧ܋�}�Qi��@�u퍸��k�o_�^Z�
S�-^��#�E�	����;*D��CX��4�d1K ģyq��86mߍ�>$2,^�G�F�M �#�]�G���9:�3HfK3��/%�k^7�9��Y�?O��ƙ'��4� �d���߅O�s�IϰC����7Џ��!all��Wt.��l)��6�ց�8���@&�����k.� ����Oc���>�_�`�4餜b�D�l�P�����$���蔾���B�q��"u��H��Z,�1�j����hhn���Ģ����k��º�820�W�-��Zl�KA�,�p)P"P�aSց�h%Ls�:Ak�@D.��o
@J��"��/^!�N�؊S�6�s:��3 ��ӻ$'��i���9�%9a��t8}�0�Jz��	 ���V��A��C2[��1��۶�@l2���j��T��k.FK �3øzu9�\@�G���@��ӑ+�r6��og��d`)*,ՏMz�����!kR�$3��$q�;;�v��s'ٗ\|س�����$���dw �Gِ!$Ӹ�U!��B(�%E�\ Q.[����>R��,3{0rpQ�o2�Q~���z `@��h��hj[[���Ȧ!ɔ���?:Y4�uY S7��s�~h�������v��G2�A�����I���i��PE*�	$Y�,�T��y���Nl��.��'a�K����)4�?�HMsg�}H�8���|����`�3@!�`�R�9���a�+A�bIL5��ca1,
2��q�ℒ��>K$�5��X,��9)鴏4k� S�X��R[�O|�N�y���ރ6���% ���Ȧ�8�ׇ�}N�p��g2 ����"�4�M��o}Ţ���{?�ڐ`��5/������_��_q��K���Gm
��7{�t�e��D9����E��?�y47����	�7ocj׷��m45��x�;/Dj�*����aǶ����Acs3�.;�����3�:Z�����X�y&�:f�=���36do�/v�s2SJ7��8��T:��MG��#`���P��� �U��[�Ż.=��T����6u=��O ����hl�{���9�f3�mF[+w��6f.�b�z4@��a݋ϡc�^X�4��
�UD�`�`$�a�Nr�����z[��߃"idF�!�q�h|��u��8���Z�ѹG�8��`	6�؃�_x���C��P>��m~� ���؁�W����\*���v:t��y{ɔ��-p�l���O�X�Jy:��OG��{����2�9�f������^C��o1E�=rrx(P���Æd��y�����f�錰:�!2��nX ��yC��m����p���}��|���� ۷�D<��ksvS-n��4�Mh�._��\C�QV��]�@���]�ry0#@ �: @(g��_������Z�v�
QQaq����@XYy")��Djz�ҕ8�T�2%�����߹���@X�/���<��BE�X�B����E)��yE$���-�����Ϟ��d���~'��� w�1��a�i�G]��-Z��T r��Y�q�58v���G�|��LL`pb���&��%s>�Ȧ6�L�L� ]�-r���bu�uE�	�����a n���VjnB��9�D"��N���D,dc�(��ΌS�0���e֣���y���	��Rx�C�"n�c�� ǭ�#âh��Mq��E�߲p�L4D����58w��FI��cZ��Z��F����A:�PE����ή�Y�A�!�߇�{�������yL�/Z�@0�� i�u���ʕ+Q���+�`�V*��5�\ó����n�A�PR8�:',�6l�ʌ������������ǭ����V���m���錎��jlٱ�������ad$�����LY�u:O�����悸4͡�� S�D�y"�:r�r�Qs�`�H�U���\�k.�+�����s�ѾRw�,������Jf����}�)Y�m-�={6ZZ�p�g�P�������l��ʵ�����݅���$J^|gvP���5ҁ���4/�  �r�BQ,^~6BU���p�*o]��eJL�ى��2*�ѫ*�#TF�q�򳤇��[�s/���w���	���/�@vs��kE�R��s�"�Vɞ��;t��q����@ȩ��� w(z	r������1 � ӄ�����Z8��ckNZZ�G�y'��'�V�Al��Xh�(X����X��h����&sE��x�\��ڒe sg��Ν�148ʁ��Zp�-W��B�+;�+�-�?��{yC�F�@~�Iy������mr���I�v�^�wOo����,r�$t 4�o�Dt7XT)�#�����\e��,�R:�� ?K�3s�K�ii~X;��:1cG��MЋҖ�ƣ���nuc=��J�MƑ�P$�� Qt��HC�3�^�t��=����f�6�#Obbt�lÕ�_�hC�~�EĳY�TY�bؐt�C�(�9K��LN�֒�.*���}����p���L�hjmBMs3���4�	
O��ȑN ���!!����<
e���j�\$Ƈ�c��(Á��:Q5dqlE~��~�NYԥ��L��bd2 0�T�N_Ԏ�o�n���$P�<�J����ѣرm;**#,@���aD�qqAt����<���q��!aF����arׅ�h���l�*��s����:)[�ӹ�9��)��'g0U�:/���� ��s���sϓ>����{5UULU��kq�W���D,���v�=��]�X���F]�,L$�(��':�TN�x�	 �D̅NaZ�[6+0�Y>G�Ё�S�f�X[�Ym��	j8��xl
N�	}�\�FGG�%�'���'e��[�x�UEF(���(�� ��Ȱ�%�sW����� M��b�
/[3��RΝ=�>�u����)�n�P��x��a�U\h��.����ڌ��f�(��ǚ�f|��������b����� G�H���>I�4t��ТU(<(����hC� �Nl	p��2J�ۓ�o��1����S�c(ǇX\��!n�ۦL���j���(i5DKx���&H�	0�
@���xo�`��q��C�$ �8�m��4�cάYصsFG'�d��p��h�[@jﺨ����y]^������+o�oy��?� �^@ك��{�����N3 !]��,!�4n�^1! "
Vz8�_,�����ϲ��; �az�֒f���M��c��[B�*��Xӊh9D���oUF��v�A2��X,δ/����8;`� ��C����^�)�kun��0o�l�FGp���a\��˦��믱]��ܒRY�]n ����.��P%q<��8���cD}v�2I/���;�E�������غu<���e�M�$K�2��޸K���W��{�]U�#�l-0��
��((���3Ǚq~u=����QQ\X�eh������������"3ֻ����~ߍ̪n�"�����Ȉ{�����>K���k��_�Ү�H���Qe��ܓ�.@����6P����]�d���8I��Q�$,R��}8��0-��H%���M��y�׍��߅���f�"@��C�CM�ųg���w�}��F��S���g�@����{���6H�bL@A0A������Y)�c�s���5�gKՊ�61s#�e�ߕ��������w�ټE��jb��k�>��O`�����ª5��#o�	�]�2X�_��c'qvj���3ߋ��8*U�U��NR�g",,�˱`�P]<��_A�Iu�XEOB$9�l��f��1��6�s&V����L�S��VgN��)R����"s��A���E��k�T*�Q�ahp@hX�A����uo6=	Fl��z�1�ǵ�7�Goo�����V��m��&Ө����"62�[�I�9�=@)�矴���}pxH���_K�]����Ӈgw����"j-l���m��]jU��	@��f�����L@h�й�HCA�(5 ��ȿJw�.���4�g駨 Q6\����._a�����a�}8�:�]<-R9Hj����P�z޽��\��^%B7����n�i���ԉQ�G.]��ݺU4 ����-�6�5w�c��?�Հ|���ݷ��Z���.�&ݽ�^��G�&�;�w3��<��4�NU����r�a3\S8-��N'�NK�v��ؒ�N��Y���t��]

$٘��J¬(\�'��L`�xZ�
m�6�m!E��2��p�V�B��EՉo'B�r�,TL' ��/������q��COo/n��Z�¥�����7�sSQo6T؉�B��� B����UQC��|y�� �I�R'],&S ��]���c�Y!����Zl���D�����-O(R���Ev7��dE���t[��� aW:Mij���)��(TOm��S��i���`���t검��|)��T����Mk�7+(\)���S@3�4�B���P\�֭[���a�]�
��߻Wr2y����7'2�`��+��ɋ`�L B��/���-����������\Ah?|�x-n��e"�& ���������/?���ڲ-Ͱs�%,Vj )h�Xd
fbal��.4D#��4�r)��b D(��/`� ��J_��à��L`ۉ ��UC�U�j��G+��Q�Q�Ve=x�KnC=������nU�����?h�K�R����,,�1"�1d�m8�	��8J�$Zb1������{Q$���A�~'�c�2��fe;��+��Dx>�U�I��oD�qiv~���[n�\���i�X �-�P&��a�K9���K�t:Դ@ �L����Hq�����pu��2�q%k�ͮ m?0��+�7�i�:��'��״��Ңk !� *#H�B+(Xꆢ5'�����?)Xr繂�%n�<iۉL@8�ڷ� .O�#�fp˶�x��bM�@�9�[C}��J�e��z�O������w�D��Ԑ.2�/�y��y�TC@g2H�"�JV\�dD�&')�A�K�K�!�����i7��]b�[�FD��Y�Q?Ѧ@��ԎH1�� �."�|����32�f;�ϩ;��	��O*.�� $d ��m"���P�X*ʄ���NG+���{��a@[�U��0�?WQ��F��y�.���>�F��SǑ�!;2(�]M:�,���b�M"Z��zH)!�rA0%�[ӹ( ���k����Ғ�
h������~W~&�r�X���+RL�y�����j��zF��KG�:���f�N=�˗ΡU[oO�Q�u~ck��5�y�pS�KuO=�I��%��`��ekLcC���f����e!Ţ��&�g���E�B���ԣB��D�B�S�������z�p��Q���MM���E�Q��\X\D��@�r��rO?���-S��� ;�G����︪ �0 ����GgW�9��ҜaeJ��K�i��=�
y�7m���a�]����z\tO�hF���;���[P�#�mMCS�g�6�h��J�\gq�b>	����a�0MG�B�E �!�sШU���2�G_Z�yr�I�����A�˿	 	th,��I����0֬_�s�pajM?�5���b���S�� ����� 74���
M��Њb��!,�S ��k����|�Ԅ����I�v�J����<Հ��Ή.��vgj˰RE5e�N}���O6�<�n~���Z�1Qe�!�^T�FQTeґ�[q���(=��A����i� �ͫ�F11:�Ç��P����7���~���1`6f�{n��P�
����
t/�opế�ݹG�\Lf���#����8% ���K3Y�ʲHT�l�ũ)',d�ݏI5`ͣ(&���"�Ew��Xz���I4�lKv� I�	f��LZӪ��]È�'Մ�(�	�2`A�y����!�F[ܩ�o"4'�T���!\Hq��6VmK%X�u� \4a;�Hd�H�Gw(Z
�S�
�-,!�֐4�e�L)8���|�eEHe�B�ҵ[�B�P���	��P�e��6J���\E�W�o�B    IDATf���[�xL������sm7�@�VdM�r	��229��{�p�(���aIW;�}ѰT��Y�#��j~����p�	��\tq��u��]3'�-�Em��2>>�[o�	;w�@Ÿ4sY�˟|�I��U�@��Y6��"d��@�!���R�~��HI�ྐ�Ӡ�+i+v�p(N\�Pi[b)�Y�eL��ϼ[���.�b���RL���s�˴@B�\[���mף�og��~�jR��&���e8~��FV���'-�A}�$�U�Q��,�Ls�U��ڢ�0=�^�"kqq��S�c��Il�rJ9}��XZ�����m���P�93c�1%�@����̅���*��4R 	:T6�ΧG4�LI?�;V��;�VS}R&��(���1	������!ȣ�X��I0������}Բ�?#ã�<;' �b�b�����<L6�M��hzvxq�')1�HiE2�t& ���J����b�d����H�d�?~� ��"@�u�����re����˘G0�ע�<y`3��r�V� F9궤�U�iK�t��	��� �w;e��e�ci�L��`��:$"j}6N��g~���d U�I�ߝe@w��E+� ߢ��~�KcNO�w H��Z9<�����	 !�$f��T������Kj�+��b�����`ځ����_��S4�����v���L`��Lq�eR!�Q,6Ԥ��z@����8���tCY��#K "�N� ��Sƚ�����`f�r�&UE
�(�|�,�?[�M�̌r��]pI���8_��sVva#WP��~ �\��h���O�X�ѲӫTѮ5 ���D�U�h1��\t&��� ȞQs�FdX,2m�֛��"I��{P�-��*��r!/����w��/<��'O�i'Xh{%�ʹ��d��$��r�-� �[2�`���ظi#J��Pp�8��7UFD����X0�P�S�TT�)v���DC�fi�Ʃ��i��Q��G�ȏD��f9ͩ=%�˽V�M7״0;}I�%/ h����*g������i���d�W@>'����	�*E@������� ����~�LTE;A�L1���+y7B�i�*���͎
�$��IZ�!k��8��R� �[�����S�/���k��M�:#�:�x�XbY�
^��j&h���B�-C�5�x��ED!=�
�i�F�W��e��XrP���q\��>���и��!ן��l�/q��c&���PʣmY�����%KO`�"�C�M�w��z�\��*����˱T����י~�ާ��⳶�x��ǂ&��JM�$�΢�댠V�#��r�L'ez����T�W<=���Ё���Ҙ����a����	H��B��j��y�[��'����w���P/�G{w+�W�{�|��&}�V����dn��&B���������$di�]�)􃘅��9]Xv�j�i�B��U��"t��D�(\���u��E��)�p&iK����t�b�D@�"�Wf������:��y�Y1'�şY��`E+ַ�P�p%��g���NIع4�m%sKvk'+�?
CĴڥ&�t n7A�<�,$�8Vu,�K�8n����5�vl�|_�ъJ���Û� ͖~o�����*���4�&iqbR�)N�Fv��k&Qm�Q�6���*�H5�]@���
٭vm����X�x	�x��J�<��T��v�aФ3�τK�U �ZI��s�6��޴�kO
�>��]pI�ۖ��D�|
���k�m�E;�j=�I\�䘩�I�'�\������7X���k_(P͸9dm}�^���ĉ�bavN�iǀ�O��"U.�e���qR �3o�$k�&�"�2�q#_���Ք��ni@"No\�`��c1�P��*���˪إ��b��s� ��?%اյJkf���M�#��Nm&�}Kjmj�L[�(�:=�C��q�hR?$�e�,t�!}B�ʠ���\Дs�L^��d+#vHEһJ �9�J�����f\�V��N)X�.��$��g굠��R���_�v��+' ���j�L!	��)����E���VK��aй.C3�@�I���>[l�c�*'�2�cN�]Z�B��\��t�~��V
(�z���D�����t
&@&Q���U�c�HG#Nk������� ���(��x�] ��{Zw?���] �R?�����������م��#��- d��K��3ϋ$2\@(ޖ�=�&��� DQ��'ƒ�5�`��<ٵ� ]Y�h;ZJ�.�亃'��~Sx"�Ԥ~����^{�K�9��J��B�r$�M-�m"qX$��I����WS��4��;�LwWE���p�ㄴ��,U��J��L$t�#�M�SŕHV��¤��B�2a�Cd�T�,��&�Y�GR��p;CM XP�2(�?) )�G	������ȻY3	�HP�����y�,��}���=�jv���������M7]�5C�x�s��ܩ3(���B)a�>�=���p�]}�XM���E�����w��p�DY�t�}�n�>%œ�J�-yo�o����j�k|���K挞r�★��b��1�>%�2W.�8e�E�~��m8�� �gfe�d��I,��H��5��ee�l:�Q�C�p�x-A���"QmC�q>�!R7��@��>��<5VԔ-�$K+��� C5U�:�󁟬ܗ�9'~n�vN��j"���/hd1!�븟t!���%N�J�<��L�857��C�/���Љ����OxH#�/��f�kE��y~��p'&p۽/�3G�w1Q %Q�	b�-�>����V�%�2���n�i���Yڹ�kQ���{�d�0|���@�Ϧ'�,���.�� �aGJ-U':������$jP'@d}%�Uw��[6;Ȧ��}�R*��j�W��㊂u��a,�D*�x��ߌ��E��y|��wtk�o���f�K+нx���vw_���}�R Ҥ���/,��O��SK@|�	��YE�����bЀ�2@R�@�P0�\�T)�II;�m��Pju�l�R��Ew_����T)�� H��2-\�q(Z,��B�#�����y��������C[�(?^]��Iw$A�<�}C�nqۍf )�A��)�}�I��̊�4)n\C���08�-e��}�}��</D�PE�Zߚ�M�$\	�\W�V)ΦК��I�vőA��2�,f���;�b$&��^�m�!g;�p��|�r	��L����8��[���*'OK���r��=U���B�`�Ă�m؝�R�� �@kV�v���aH
��6�Y(Bi���������J�{�v�k̮�h�Y��ΰ��8g�����6)G�(����`�܇�o������Q�/�� >��{M��l�g�^�,<MS���R}�puexE��:7�R���+�?Q � @��$���s����}]I*�^����C��bڶ�@V�V�-�&ͭ�!�-E�kLl�S ��Y� y��N�﫽R�ᮀ��y<�:�4�6Aq��N���G[�$A��8�n��Ο�HM ��
���y��@W����&����'W�CS���4 r����h����Fx>�IK(���e�o�i�!�=�'����i(�����hcn6�3+�LK�Ci����_�O������Q�`-.��d����~�GpӺ�S] �O>Q�/���^�. ��X�N�J��B�J���|�Cx���P�|�0���|`؞�z�h'��"���P-T��t�����-uy��vK�>�>�E��l$�Pf�H�m���'�-�:R�� �>�ٝ�x����G��I�q�2	H�|�S+������,`���ЊpD����<�J���:B&<{!�H���|�gVh(����B[baA�P*bb�:؅�L]��0GKY��<x��@�!v�����DaK���=�|�N�(z
�E�� Zu	2$���r��!�B�q1T@�vq�g`
A��,��M۶��Ϡr���~�A�L@�g�p5�1�	��,<JH��0Yp����[̸ ˆpRu�9�J��;�rZ�jS ��W�)�ļ� R��m#��$8%D�nq��-1b�Q��|� <��:9��p��x�_D�f���$h�1̬+�ũ���:$�!���Ԝ��������C%��ܾ�KSe�^hy2�ιP��X�\XXU�.c��q�hS��b��PO��h|8�:j%��'jc	�~q��R��SP
��Q4-�-��	�/�@���h��E�̩�x�� 6�*�B�Ek}���(J���(�9���9�n�\�����ɹ��
^��"���ϋ�t��9���wln��`�Ǘ��fu٬�=���D2^�M�M�S�0f����n��Aw:�E�5q�jgF� �,���)�_j�A �����}�%^.zj���E B��`���Vm��M��&~�?���K���{���P�
����
t/�opế�ݹ ��0��Y�ۃ��-|䑽@"#'y,���R<-,zB$1'!��@�ź�*��t&�R��A��
P.�(� ke�gR���3SKO:�,��"���C�6Ѩ���\xQ�z+��q�A{IF�`���:�>����F>+P�G(�u[D���f�.l�]Q{�W��#��dw��	oih�}�}x%��?ߋS�t#߱P�A ����$FW��J�Ք�	
ƙ�Q��V�T� �5R��J�s�9-��NM��J���w�X���Z�u�x��aJv@Q�H�H���U��X��`��i���;�����{��ƪ�!,]��	����P���!l�I���BL����3O����)[(2eH���d&�U�*��	�:���W|��S
j�*�P���Q"I�t�"����-��I
��7_��k6a�SO��XQT�,��$E�����O��f6�
��T#-�5�PA,��BO:� �J��"@�0��+���$��p5mS�=��Z)0�B:յ�����tO
p�p݄���/�����'�0�N��c�׷c����Zжz}��& ��Gl��K=���V6�
Dp-t�^�Qu�v$�E��qrV,��+!�f����礖�lZK�{O/^c+k�x�y�R��"�|ҫ�%T?������t��6F���� ��^�q��]O�����C6^#��-Qm4U��qƖɇ�4��2�w "�0�������BLmxe��IPѓ��,�lӐ���~ �e` o��x֗-�~�� ߝ�@w��+� ߊU�~�Kf�?) ���&�VA ��~q�^�"H\�}|g��F��-�EBwγvn�B9j�/��"���P���ˣ'g"�:�$
����)�'@������K�s��ڊ1_m���`ٴ�d22�;�E����-m$�N�JS\�X��n��a��%\-KuUA��#��8�"̍)�ۍ&�b_&0�k+��ҝ�E&�A�![��-R~�s������)�<��q4�^���B8��(]!�2B)�k���6�^�"8��*�|.`���~�V�z,6�H�c�t�k��Q���!l^�珝��'�Aqp�zC47���>�r�N|���k&�p�fO�Fmf�\Q�R:�;�3h "T��)J:|Q%ا�������D���uhJ)Mg�S��ϐ���e&ҊN�N�Z��6)oM`	��ad{�"�'=��؃�lƳ�?�Ve���A�&:�C�
�)q��JM :���7�  ����C�u�������{��a�.���^�c���#�'MML��d��&]J����ƭ�OH�y�rZ��^��+�t�.����
��"U,�$�e�d��'�y_���I������
�*�Iהۭ�gR����32����eDj�2�UT;���FЬ�+����_!���xzʥ�����>tF����0�׋K���^�E�f.NA��M[TS�ɢ�
��S ��~_S��0�^��t�љl���Zw���RT,κ�����	l##�c�����#�6П�����Q��1�o��;�"���ý���q+� �q���A��  �T����؀�881��Gُ3�1]����C�+����Ti�/>�]Zu��*
n��A�.z��y#DO�B@+V��޼��T;W$[M�G�)`z����	)xۉ�V`�Ĺy,6Bԃ�F� ��aRk�\/N>�"gq�)��@���{+b�X�hλ$���Z��ҝ�&&�'-���bfB]03Q��`��Ț�X�"�=Y�&Wa`l��|��8��A���O��9�7(m۪�?��0'+\sҠ(��Wv` ��m�5�P4tEya�\�h�}������;�}�~�)T/�
��gbo~��3���?|�lۂ�{�b��a�y�L�fD�c�i ���!8PD)yΰ����V*?�f&�@��#Š�1J�QU��i��Sp/��ӿ��W��U��4)�ȠP���� -&�'Fz{qӶ���#_@s� Dm*9�i�P�XtS�����r
�q�l�.�;baҦ4�j���֯"*g��|)��Qb�L[w��qkY�$�6Y#��)��р���) Q4��[1AI��" ����X��"�qaPa��O�S�О�fb���êd<mɫ����dMe|�^���;�4��)Ǖ��b`��(�����:� �xF�j.�t15��Ӌ+ ����I��+�2 ѧr:�J��쵩}"m��[���Ȯ'���`��É�g�mlޱ�����i���ޥ��h;��YiU8�I@�l�t��s��ȹ��/�0]SK�9LRԖ�i
@,(
֚�q�߷O4 �B������	l��依�vk�o����/��^</�����o�
P�^m�B� ���C �G����xqqB�v[4�>Ww���Ja�jZ[��vqk6<��(a��l�
�h`��b�'��7mG��m�e�j$JFeiu���|���ũ9 M/D&���ǒ��$8q����<�Za�(a�k(N)Xb jIq+Mhv�ydy)�X�����Au�31;kx�@,fZM�G	�3\D��ӿC�!u��	�T+F|��3@nd��נ��X�֤XjGl3~hp��R�Yd�eHrG�qfb��6ږj�&Ε�Y�
vOg/]Bl��0�CД�y2�җ�En���o��֮Gma���O`t�j�x�-��ǳ{�����qݳ���oU��	4Dߡ��2W	�%�Z�I[D��R�dm��o��.2E���>�y��UT��+z����j'gB���o�]a!�ƦrV�d4�0:,6�� ���M۶᫏<��ܼ�nZ�*Q=�,v�;)ԉL�R*OGd�6X�*DCa��J��q �i�.z�QZ��1��N���'��`K}J_������7��.5:�}M�T�G��Q�~�D�3h�1��6���ά�(���0�lنz�.���m�KNܨ]�� �x�&HAR���c���@Q���j'<}N�u�#)��ّ�9<��T�g��,�Y����^g*��Ҧ(�N��Z/�S������j ��4m]4l���L��X�)��۷c��Y<�7��s$��������O�F��@��H���92B�#��mf����z:P
F����6ŕ ��C�7�a� ���8x� ��K�as>~��~7��C�t���e�������
t/��C��ѯgv>���']�����������{p��o[b��b�E_&p$x���u�ρ�\����H����(%�kc�x�=�l�@o�]�+`%�_o��=�=���W7/]�S'��ĩ38z�Μ�A���T�gP�S�g��2Pk�h���t
ºb����C��,O_ہ����P�4�9!i�(�U�h_|��@�f�S.T�ST/|}ڴ�hSo��+������ʣÀ�bnnNB��p�J�ݮ�v@w����8�
� �PDЪ fQb��f1�z�$��I�VK���e[��Xg&�␓ժ#_(��19��G�    IDAT
G�?&�#��8w�,Ξ>���!L�����1}�6�E�f8����3G%#�h�D�7Y�[g��y�MX�$6�⢦��Q �>K���c)�Rw%vn١��	�v��Y
�ڤ��m��^.�aX�0@���o1�BO	��"Z�/�616��^�/}�a,-,��̂]��T���w��bQ�4/��-V�5;Ԥ%i �*}�i�mR�T7>d���K� C�_��r|�������g�&>��I�pEd,R�����^��W�ν��(WV�eZ���HN8����C;�l6� ���ۋm� a����"�\A�q��Q+������8�^������e+`R'�X!gLW���S,F�~r���3_��U����
 T���W�x\1�ֿWL<:NoiA��H�7��w��l�cdsY�����������'G����M`i��E3���]=v�{�
Q��C���Sv�b�!۫�hW����vZ��|,S�R ��W��m��{�a��cr|�@�фk�*��ş}+V9��%�j�M���y�v_�]�Y����=-�+�b�s0��TRy�6�v
�{�2>��n�^�d��{��6�~�Ba�D4�{Vv��sbl��j�ƚ���~�Fm�@r��!�]>�jmA(I��#��,lD ʢ�Bcq,�ʥR	�r֮߀��1X�����><����s��l"��Zdcf���j��z^`!�X�qGc8��v�I��TA���*�-�%7#c�trr�NjqR� �kW��,�M�t#��mN.��S�$
�;6��U�0�9\^\Du����$��=Q�	3b��Ӻ�Uai@���me\�t�) C�h����88�s��B���u��1��`UeĎ��XYRXh��;,�=��R�b��@����D�i�5��gB��?�C��`�,�����R��P_B�X�إp�Iۜ�H����Nf�R��>'%����`U���+tF�ʄA��  ����a��� D�|�}�X�T�y�f�z����?���s"�$��4%�*dm��7�W�3##Ų��9�1N���,�@��z��	IQ/�uDg�U�j�8���	��kҴ�����!p0a�y|}�o\�͆�INʠNV�A���?m{����4�����������4j59w3����,0��B��$O����`P#�Rj�4�ף� r�P�%�/�A�ʶ�?S��*{����jFĲY����R	F_/B�rd�[�Pf_}�O��\�+@��c�%���tD4��DS�3W��k�l"�ω=�L��(|x�oy��q��s8}��2�0¹��Q,�ɺUi�M��
yn�>��)��b1/��C�,� LƏZ� ��]):�����099)S��{���T�ݎ1V��߾�_�=�h.��;��n�]�ot� �]���}W��{	 ���f��>�xt?�N�ж��Im����9
,���b"՗П�b�D	�Fcܴq���6l�v���KN.�:����kUa8�LM섉��$-�{ͬ��yA�&R���O�G�b�������ј��}��Cp�C�4�N_\�|�6�S��ER�(0� Q/�"�˳ܱ`r�X ��EmED����)�}��S��K�COg/�Pኑ��ڐ�:!ܘC�6�*��j�鳛�A��0�H��-j2%6�CeI��%���'q�HG8�TŶ�+�
�j�kI�:�U!�ݔ�ob�:�F�������t$St:�D��'�������Q��P?V��{Q;{�>���%D�
&0b�cHǗ6���)��.
�.��:t�q[�-�ʒ��T6va��t�0B���=��1)�i����U�K���<��Z#!9$,�ʍ�o�)��-�xe�Z�&���P��T�7�&��Ve�[����,����a�bnf��ً��^�\�C�h�<4"4�F��b��T^Mȱ��G$)BO��q*��SC�6��)u�b�� �e ����૤{��� �[@�ӥv&F>k��8�R9�h#�ϣU�q(�M�?��"cȴ��R�Q�
(+�(��h5�������
 �Z>�9�˙�y���TE/;�4���ߓ���ZU 1�ΆA���9���F���T�j�*A��A.���2��J+���P�͒2E�a
3IlX٢6��~Ѣ�4��P)��~$�� �LAt8��T� -����꛹L�t�~���ʒa�tD��z�e]	�5WQ�x.
���6}�y�9,V����|��bh�mwS�]y�Ա+�]��4�L������9��B��lL( ��l�Z�J ���{���  d���_~�;19`�]�ūw�ܭ��++��N}+V�{�|+V��/�  �{�b�@4�p�ԑ3�Ҿs8t~~B�;]oҔov�]t
"�'�0֛�X��XO�7ܻ�_7�M�è\<�'���/9��jt�F�I�<��/��^�d�S���G1\�F���S�a���X{���S��=�����Dyd"��Ŧ������)4v�U���������Em1;O;i26"�XHq���	���v$�W��k
ݟX���R��"x*�`b�5�s��]X��6��R�.�k�P$�	�� 	ʩ��КX�+Q7�Y�NN�mY�����ߏHh>�ʧ
"�e=�0��6�� n@��1�ޖ8��yl��S��دc���LL��/������-(ZS���rB�B��C�L�@�U �p��l�X,I�ڬS|=M��h�Y:�q����8��;�Lێb���Kڽ�W�n�l�@Шr��%�B�pm 2166�w���X�v��&��M`jj��'�W�
��]������
%�z�(}N�&y,nNM?"#�5���5UF,�4��V�B�Ra���L@Xk�����05I����+`av
y�	�)���?�O��K�;�W(�$k�Ǖ���߮��e�b�Q�,׶���礩Zo!�+����(|�N#B!����@u	��>Y�|>�z��&�ٱȉ@�gI��)r�G�����#��� 'qKKKr�Rw�y{��oqn	����S5�6=�sYXԁ0�>u�ҁ�2�H��8Q�y</@::��ڴbb�\�:@dE���� ?�[�d� ����(��e�cۮ:ŵ��-N`u����b��)+���¯6?Џ�N�sU�#�W^c) ]�e�3 �����DI}����n��y�w7�;m��w��nϷuH�" ����-�x����u��}�g0��*|�1�"#\�l;B&h�7�`�x=v׮)���ȴ.�~��؏�k�� @�!�PY$8gJw���E�3�\;#EQ^�<��S����Gw'`ÖM�f�u�{����?��\Naf~T�X��Ρ�h��E����B�(C�]��X�S�s�"�/UE>�N�B֔�E�믺�r�P����$Hjzv�m�2JCÒbܤ���KNv;D���6��vA)��T,��64ښ�N2|����1:1
'�����8��P:��@KΡ&<��\��
�PgcX&2&����wEfd�����3h���d� �=�4��Y%,6������wD6GO0N.��^>�d=8�"0#Шךr�)&^�_��v�*�E��4k��,j%łt%���	�̨�-��5�����eJ�q�Zlټ������03sYޏ9�qEkԎ<�u����?����x��_�]���� ĉ�g�Ȍ��	�!ŭA�T��b?M��G&��9D>�yYmG��*1pS��UY)w& �FY�UM�H$]�E$���Iiòc���"lT0u�(J���V��FN�V 9�<���h5�ͺ m%
�׮]-�?�>r���RU�]ӂ�Ш5Q,chl�Ob"W(�V�ņ�cx�}�೟�4.�;#�9O�&	3-9��t��LB����X�rY�������ai~Q �b�"�8_K���,�-"?8�-�n���GN��<��	%�/{tD �x&)Q��� %�N��Q rŝ��Rҗ@���
M**��T��r'�)/��1�P�S�9ok�O��%��̟e���̥Niڕ-��i��& )%�c���=I)X��y����9����$��L��
���ۺ5Է������
t/�����n�7}8i��|re����s���g�pq�Ϗ��;�Ќ�#��sc�ɣǮb�d�޺?p�M8��1?xP���R������+�	Q�.��Ϳ��g��eЙ�׵Q�.�B֥���bu�0@�܏�������>�S���L ��aj���R�^�A�ɣMw,a� �]s��V7D��j�VC�E:��t	���)Fv���BI�YNo}##0ry��W���&Ü�8B�������ZO�7mS����B۱v�c$"p�(��T�#�Ϣ�jH�y���EA�][�$� (0=���'I�Л�-2�u�$m��J8B�51X.c��0�ڋ�\E��m7����q*�����Y)R�6]�B��U�
9d�9T�0:1!.jqxL+�2����nf�$��4im!��C�9���A�wۮ��j�엂U�;�*֯[�{�؁�b����ͧZ�	��!y�6��+^~7>�k�vų��}��������7�s����}������5�2u�o��3l����|�BZ�ur*�&���qɱ��|����*��b���N�H#2u8���c}hU�`'tw
PȻ�^�$6�>��&����!�T��B5۹�V�׍ڝ�G��Ѩ��t�2.\��V3����`���x���1sqZ&N���[o��y���ڸp�4���#��`��ŋ�Y�yJ�mb�����@oo������78�\6������*�ǘ���k�䙳x�ˏ����wݏY��s>��؀��0|�uጎ����d4�$Dp�D�� m��E�וb�o�/��%O1%R��%ۇ ��D#�NE��o�UP)�>�lҰ"��o�Bi󃎳�
 "�Lm�Ѩh��(Z+H�O$7� ��s@R R�2�q�ޟy�L@젊���u���?��o�=�] �=s��;������K��*(ۦ�������8v��J��ah�w`QF���a;��ĶUy\����޳e��O�՟��JYA���J4�ɢ���%TjMI�.{�&%@[r��XZ�J#�Q�fPt-��a������R� ���?��u����'~S�!��8q�<\^�P�-��d\�`�DC,)�U%u�B]��)݄z�	,�$���!���dD��~m���׃��q���D�153+zǰa�m��E��:2:CrT���fI���0Q��-br�(��Ě���9�jgI1j5UG�k*��� �u%�<�m7%���-�) �Y~���S�O�b����DO?�x������0Xk$���11:���Ʊ��P�e�7������BO:�gN�����P�7�s��w��anfF:���I��	�;4'8a
_��W0==#6��b?�U���pe��b:��������4��,�=2Q�C��R����b��Ԧ��&.���؉��˿��/�`;Y����ؾ}^v��b�R�������p����#����x��g�]�2j��BU�*q��LX'(����҈��[�d2dQ�`��Q�q�f��^���~�A[W��<�;��9sN�����qa� MNo���>���Yр�˱3�����OI�x�	<���x��Q��U����*|�_Ʃ����[�f��zu�x�;�n�ۖP�Uk�G��J��O��gwcr9��E����Y��x�vD;�믻���q󦍝}8=3���G>�_���F�8�e��>�ܡSp�=8�e�����9a�|�h�* �bk "s6�TS���x%@I����^�ke`�k͉�o13H2z�4��gm�H�Y��*u$�$dv��%S.w�|Q�&����% �˗h���r�����v��t�� D\�}]� 29:���>�z�����?� ]���T��/�] �=3�+�b���"ġ�V؆o�x��i|~�I���$��#+ �<��(e"8�Y��շ�����a���1}���ۋ�p�U��Y7�¶���c�M���~}��g@ �K�%��X\���g��s��i��f����b�����Y��M���k����⣟A~h5������������J����~C���O�wn��!(^�Iҩm)��XO
 ���E]2])Ö;����(J��h�Cp�T�UQ��U���-��q��\��ŧ-�Ov�M��P�o2G$B�X��rb����c��P�Po6$��]��F̉��,���Hr%Ć�-�ձ�U�$�
\��O� I�1i]Q ��.F{p��!�զX�2�:��r�Z�%�]5���݀^y7�9a��k�S����MΜ;���LMM��k��]w܁�g�J:�*�ڢ��+�h��#@�]��NJR���![(cna^+�R�*Z�g4 ��em��5kU��֭���������{�m�,�'��q�v�-ۍ�{w%���!�fg�G�Waǎ�q�l]=�yn����>���>�/?�$ⶍ�O?�n�~+F��_A�I�T�:i���U�d�I��� "2�2eQ+�sj�ڸi��v�Z�v�V��\����_�<{��	A,?��s�P���˗q��>�N_B>��������w����G��#�N?!b�k7 n���=���G>��m���lܸ^� �p�x�Mx��`�ރ8�".NMc���Q,�E#B ���d�YoyX�v������x�~����~�_���*��;^�Z8��	$l �ʶ���sp�4 ���Z��	kT*��<��9+��i.���z�D�`I��+%J��l�+�N��X�?�؂��P�p�|�h��P�V %�[�	X҈�E' ��@2:���HZ�.�c
 Y�j��cس���h@8I)Xh������P�
����
t/�opế�ݹ���H��@
��vO:�O=yg"�3� 3�ϗL3N���sx׏܋�����e\8���z�#h1�;��k�BAB~xAx����r����u��N&����И�����
.r�����=���}k�����q�ހ(S��xl�sh����TpӋ1f�#���^�Da t'�VQ4�"�%�����N��Xx��'e)��� ꈙ�a�X��x�6./U	zzzP[�!�ڈ�f�B�����TǓ�w�&PN�5�[F�Dجe��ۃ��IԂD��@��
���rg$�?$tQ�v.�ЫxJ�\���N�#�f����E=��hT��>�LkG'p|�U���1Â�2ݘ�V�V���7`�7�գC�~��+��'>�dvv'N�PE��7�PZ��#\�ӧOcaaw4�c8��-W�h[:'jO�ͼ�t-�a���/���cݚ�����F��Z��_��_���0�zꉄ���n��n��'����o ��~��rL����+��?���#~�>����܉�{����kb�Ru� v�"v�t@� �h�a��k'-�;q�bN�X4�&�tsm�|��7oƭ��b���1><��,Oһ�3O�MRgf.avaVhM뜀�iM4VY6n�s������]q�:~�yT��K���K,V�bO�˺p���2q\[�#�^lܴXO� �|Q(�7�t�hg��Z��s�A�B��!��y;��^�~�r��~�/�_����.v�y?Z��g��I:"�X��m�Zi"?9����^6���4�<�I��4�t��?��G�����@�jӤ�+�L":A�W�48�Ny)�����&��0PQ8uJ�ƧӒ��X�v-���<.��lG:G�
���������N�l��5Մ��#�x	@V��c��]��R�-р��5ғ Z��7����������Uw��+нx��k�}��  �E,�����<y�4>�����v�h�%%n"-aC���������m��W���c#g�b�tV)��v����q�o�g_���xR��Be��Ρ� �׌�٪�#�/���,�����G��gv,�v    IDAT��K@a�݇�
�%e<|�A6ʁ�S�Uw�D�{'A3�j+\_��8l�غTt07}
?��?����DO*X��q�RA����>\�<-��'����#��͖`y��֧�0;�tS�l�(@_� �b���Wt�+������;P�4?�J���m`�����d��W��$@��4[#J���5[��A�G)����
q���r?�H��e6��"Tڴ*�{������GQ��'c"��h!��tkx�ݷ��ඛ��uw^�����ɞ����T�}��l[,NYP]�4�?�П���)�r'����,��,��l^i]t����T$��C�z�����z����?������=_:��f.���o�+��p k׬���8z�e�t���>�������_x_��c���ް��]@�s�)�:^�*��,��"R�l�i3�]c7'�i$V˜xi篶���s.Jyf�Ě��o�u��_~�?z=�է��{w	H<?u~ܦ�_�
L���t��䇾���g/!Z�uT��[T��B[[j��?$ǉv�V�0�ľL���C�� �ib`��oc�֊�@6_�m��0�< ٷo.\���a�R��Y�a�P�������
���?��䃿����418��U�٩@?0lP�3nŉQ�h2A@%b�,J���+]�w���D'��v��=^kG:��"F�����T��f�a(�j��S���ӯ ����a���{�W�B��\=Q@WA_Wj@H�d#�v�k֬�$��{��1��D& ����IH\���z��n�E���tW���
�����[�}��
|�W`��@L:M�	���ϝ�?<}3Mr`NH��p�N�c]��{������5��⇒Ӈ���@/���!�qQ��Glh$&n���0���uלڕ$�js���?������.Z��t\�{�Y���7����_��E}�[pf���Vg�Z�1�At�Ðv��h�]�P��J(0$lQ �0����c릵x߿���U/�|��$��r2����a��gw'����v�l�l�ͥ:�h4�70a�C\�����}v�v�LZƑ�K��UeY���	]���e���ډ�v3�}�ǟ���'.�e�Em��瑵ۨΜ�����+�^�z��?��<�9�B�q�B��B^F4��M���2F���p�$�_�%���h+�Z�r	q�������6���z��<λ�H�O]D�upi��"1n���V��K\����������Ū8Qٮ�Z��'8	��`�EhddD�$T�\�twjΟ?/ ̿ ��%َ�w����%3����/����_���ò�([=1)����qlٲEB ���Y<s� ��o>��pq������'ag�¶�uϜ$Y�#�-#Y#Զ\�8�V�&t:l��*��$b��XyT.�TQ97Ķcx�[^����U_s��=�,--bz��.]������0<<��=���{gϜJ�֞ה�xϯ"k���:���4
nfk�NȉF�Mϗ�J�d;@�an�r~��XXj�P���|�6nŵ�}�q�����s�.;�'mv��Qo�p�y��~���� x����� L��������>{����(��)nX��1x�@ϴw5Y ��M=��ajJ��l@VN:�*u-KuS�Ƽ�H�.&���)Z{n���k�fX\���ߋ�&S����B�ru��2�KQ��Զt�+=CVhYR:�8����	�l_lt �A6
a��
�����JH������~�Kz�E��Kzϻ�]�Y�'��K"r�M�N�����G/��}�pn1D�,�u%�e��d)��}�p�8~��;�ا>���YL���X�B�ba7_������y3���"�܃�8�;IZU<��C8{�0Z�E���Ϣ�ԋZ��b��u��Į���y���X�z��q�\U&r������Vbp�S�}���\�^�)���;��?�:���k�Cg������_L(r��A�~�l���Iq�a��s�y��l���/"N����C�+���Z�����&�����G���ɩF��TP�����N������/c�c�?����?�<��9�8�����
��8�}��*�Ə�]�/���D�!L,nAܥ�A(�"�	�fX\��Gp��QT/^�	S����#�uM��Z��v��V�}=��@B��B����)����률u]vF�x<x���p'Eh��k�f�:���N����8y�K�Q��?�z�~��8q�|�AL���[��fq]���~D(]�sH�"�}�v����J�<V�������16:!I܍Z]\�j�aشir�"N\8������o��-�m��'/ ��~�X8S�B[�4��c/X_�##c8s挘-䉽5�.l���DƠ=��4w# r�� ����=p�?
@�"�p��Y\�|I@O_� ^��W�:@?4��1'�^]B6��Q���a�8�Q�����̍�$��HhkL�P �]�`�b#�k�f�f0���ZN.+�*����>�	�/,!W(˄����'�	�{���	��_�*� ?����7�/=	+WBSC�
ڔ����0Z,�E�eJ�h�8
ca�R�xRj�w:=��j�
����j��\��u���� D��U�t��9�!���"u8<x���d��_/ ���9!�q��^2���(�?�_	h��+& ե%8I[ s@֍� ���꾾�W�@�tO��
�X
�ɭf78�[���GO���yT}�����j�,�e]?�÷�^�᧾$!�Y7S��0F�o��}&n��o�5�^8��@��=�#�w���}@�c��t�Y��/֑���u������A�]@ad��$��gq���r+�d�P��KD��JR��9=Y��e��;߆�zߛ:�q�\%ٴ��ݯ�gg�k�;���s3�;��~�U�YYI���k,��m��?�6��k�p��Z�a�t���h&�����g�;�����s�黳�%[�I%��A���^@�Q���rE�XPD�	!��MO�'��w�̙������d�x�{|�w�'��N9�w�|���%P�����:� 5��/��u��S���WQY?���L|��>���w�-�c�?Ǝ}Q\��;������i+T.�XcS��r� d_[b��l�K�j��MC��Esq��#��O_��k�����T�:݊,bld�� �$�P)?Ep�u�V�w�}|-]z$�������P���[���܏��1TTV�����q+�~���/��x�QG�w�{���K_��y��g`p�+y���/|��_�FY")#$�݇~����0s&$ŝ����0�Q�D��;4��<���M��v��#9M�ZUX`��.����%��U�q!�X���&���nϙ��K�8=\=�T3&PU����]}��=������C����������D"���Ùg�*���u������8S�1�	F:����"�\
e��4y=�u���AZ!	&׎��I.k2�f-DiU��ON<
�]� �p���k��g��E,��8���&���n�D<�W_{k74��˯�[vcOk7 �9�B3!ʐ�AH�@�Z��{!���I9��tw;
 ��w�A���A��{�R��M ����2���֏�9D�*�&g ���,ܫ}�K��ݮ�zBI������Ȃ�U"NgSS�k�i�z�`i����W��* �O�`M�S+����;R��?�ʩ��k����X�]7)��ANP���k����c	]@"A���Ǽr+���;�<��X���t&U�
���F]�,Z�B�p�?��Ɂ�N"ڏ��ط���QS�N�t��?��X��'��ϯۊ����0��w(�T��UD˰��iG@H�N�Dԉ�$��dHvfb/��3V�rǞ��μ�r�c�t<*�WH��������W7�m�9���4��|�!��?�� ���c�N�?�>�:�p�Į��3��A7E8:�:�`d��j���$�L�8	>I�ko�9��� T1�E悑F�_��O�3��̈_x��p.��SH�,��E���C&%��Ƥ��0*KK��ف���\kb���$jTS:��ƺr,[8�ƿ��vv�;�$�c�mc#����TϹ	~��shH�[շ��-�L��U�>R�*��q�:;ڜ��~
��{/���� �f?��MN�6��{���z�w}�Y�r%�~�x����Q��/~U�x��E���O� �72�H�2�|_����j~N��L����(~��?ah ��G�}�C��EBhZGUИj�x4a",%R�By�=�P��M\�a�yHSrb3l7?Ʋ] b�Q����.ƍ���m��6���!�+��ӄM�6���5�u�3k.ο�l��}�C˔�Bt1���ȝ HOW�;P�`��t����Z��Y�7�����놵;�,Q�pD/.~1�Ƣl@]���f�OQQO��/hk��uOsH��7�3��/`�X<�����4Jj���e�m�Aڔ0�  "x�p�.��a�H���� 4E*�,"'�:q�
�'�����M2
�˿����{oF^l>yrA�G�+L�h�H{�;Пt�<	�`�I"���_N�����<�+�ķ�7�q҃L�d74�&!�b�ϟ� d�������R���~�ØQ� ©��l���+0@��π��?l����$��D+>�����^ܺ�CNO�6F�\G�i8cin��5¯�s��XI{1����-Fu�̚����`q�c�#Y�v�yӫ�J�&��T
��#��-������J�+��՗�X���.m'�V�������S$�cC(�
پF�7wJ]Z՚]�Ύh��S����jiE$�����mj���/Ü*Ih�:�vdS��:�8���@q$ME&G$�������v�84�X8�V��_w;�=�<Z���Q�E�D���(/+Ɗ���^耞J@�!y�#N������=��⧐s9̊���i�O}1KB,Qc������`���@8@uy���0ѳ�ט�<
R(��N�ue�+/ƭ7]�7v����pF&��cbb�t��c9155�:�>��5H@�����?���!��ރ�ŧ�~&>|�U(+-��ի�/}	ˎ:
�������_aժU��ր�|�+d�+�}��ΓO>��wv��lhMJ�M)�!q "F>��#�=c6.�1�g{�>TVW2n��=}�k^Y��olE�%�e8��hI�D���S�#OۘC?P9�/�g�!�mB�5L����^�x}|����
@QP�h'�3���?��n��5޽��.O�wv��n�8�����6bdhӧ5`��#QUY@bq����G ����!>6���m��T8z
~�=뺌��^�P��[$p/���ÐX�U\Z�iMsQ޸H����d�Y�T��d*�����ɧ�go'�d�O�x}*JKQ[S�k��3f��_�mF<�L	�����-�Ɋ��	��\u+�%x�ي���w߻���Y_��"��/�h�',p�D�*h�
 �,�]���L�r'� ����]�|&�UE8��-�H���� >ȕ�6	@�Z�uϋ���ӛ�t���;��77_�"�+Z�`�` ��_�<�����T�JB���V��\�) �O.����[+�co�3<1ήA�(!e���a��N���&d(�Bϡؓ�i�p�	s��)�����|d�AΓ�(Bqy#/9��w�/~�w��K�����Ho֬|M��9*t���>{6��p�y߃X�n/��� ���X�>8���'9>����	ɂ�]_��B�(�⸣�����@��pK�)������7 G�_R�I�����e	z�E�v�pڙ'bQ� �����n\~�u�J�[&L3��������qGm4��
_{��/�x�Y�@	�_Ѷ�YP8;���1���Kq�+0G�=9�9򤫐�=������0j�*���w�$4Eṽ��'n��� �d�ԋ��K����npi �ա}�N����Y��ϴf��)��F]e�!���J,[Є��*���س�ii���� �K|~>UCcc=l��|7x��5x�G���a�K���*�s�����-�뮻02:��~t?�>��W�8���=��%ť��{H"�\�ҹ��o`ɒ%l�K*��q��K/��� s�ItN�.D��d?�><���OiAg�����,��X����k�?��Xj�z2�6Y!�9i%,ɓ�F�M�w�M��EY0�"�ұ	�p�^P�I2��KJA3(�����C�|p}�ܲ�����'3>h�S][��׽�������+pƩg��$Iv�J'��M�^����8�T#��#��WD.�";��	���dt(���ؔQ�Ԑ�)e>� $��`����K1Ob����=�xt��,�q��m�d�bM���}=�|¥�]��>x��j�^g�������=M吡k���r؆�UK���(@ByrsSܰJn��� �5. �4�|�8Mzx �B��nRo��O>����?|��ǒ�-\@q�A��������<��@H?# B<L)�ɮ\��y���Ɉ�8��8X�G�}��X<�a��`��y�(�`��7�J&ن7�8��uBSe Nr�����UL�Ϳp�.��bO}���+�����bn�!�l����k��`�r�ʜ�GC����ጥ՘[b`�O!��:��O��P�t$f�[�p��۱��+20���J��J���g� �c����zd\x��xj�+x���B
�a0�@���y`�Ųd_K�{E�'��3��d$��H �s
~t��c�SV�U�[�O�r��Z������I�gxx=ÄGV���8�ӦWc���h�=c���ș:��~�2�|��BKߘ3����O�}��γ�o�hƁ-�9ۃ�d�H�$+䢨,���O]�V�EWO�|�����Q�&�9����oF��jG������m�������L���]ad�,��L�����fX�8N���Ú*``�Ng����^�ڲ B~sk����wz�����zA�jC����rvV"��L�.Ń]�v�g?�OK����Ԅ��'��n��ϝU+�śo��SN9��9a=������Ȣq�7��o�3g����h�¼y�i�&�������c�g�y&�GF\��5������ׂ,H�]D�*l޾��$�`r��W׽	[�at$
Uä�-V)��-0��/P�=u�I�B��$��`B���x��(|�:�L{+��_�Q�up����x�{lժ� Ė��g��&��+�����N���I+V��cW;�mvt�`�8����Q�`b�Ff;ǓEQ08���D�8��G U�H岠Pr�����V���cP3w��{�&'���mBA�F���O<�$:��B��|�JK�81!:1�SO?��x���[���П'�}�順�Aa���fؐ#V!���m̠c��e�P�Ncy� 5*�GS(Æ@<��n�Y-ya�{���u�,�l����mq�WH�JE?/8g����b����q� ��ʼ�&���&����y�	�>t���qmymɝ��0�Z7��������f�<R�7֭���6�|n��J4U�S�8��) ��~�M���w� ȿﱟ��Y�--e h����`{�^�؁��b�����s3�X�	�p��"4�ؽ�%�ad2i�^�/�yKOE���ߵ�lp��1�	(V>���<�k�1�5��tѣB�l�q��xy}3���oa���D,�EˁQL$�����S_�U��L+2�)����.9�4|�×@��+a�ֽ��w@
A��F5��,9@6�����e��M�F6���q`�I�TT�r�7}&�}�p�"<��B�@ԙUU$�w���ر��P�t�i�3$MSɩʈ#�AUi��|
G'�浍�T� �N#����_�o�����XP~��ù���"�)Bʦ��E�)*    IDAT�%�sP�h�8�ô�jlݴ	�K2bs�SX�Ş�H؋�/µ�fv�=]��ծNawk�C�c������31{�L.�IB#9b�0�?�z{{A���_�O}�f�?��y�3����;p�E��=��!�A�=t�áb�z뭨�>����A���s�u�m_B[[���Z�r��`W.�+2�� �{~5��)��+k����{�6*.³/���dPػ���F0�~�@ ː��]\��rpC.�Q�[p�b�&ru��D���Rf��Ƣ{u��,�����>�q\s�!���69�e�Km'	ڋ��ش���D��(��3�p�y�
ۛ7:���X�q!�md3�DA61�4,�)�D����)�3��\pi��Ж�S���@�����0L˖�ʹG
�m-Ng������r���?���PV^��o��\&U�ص�%K��n6��w�����O~#�r�[�8�E����Ͷp-v]�)�V�2�`���+�t����Jr���@	����X����6K���� �¹W�aw�ɺ���m!|龾0)�����`0b>h�-���rL<@���E.�c�?r���e�̞9e�ֿ��4���|���0�B���9Ǿ;��/��wX�w�0�wX��}|����{���1����a!%*x�����{<���,'���� p��Z���*y�m��ds��o�ˎ�E�K��묧{��҈�%�|�7��B��5��<::��O>��Կ|����G�F�a )c8N��~Ds�T�U3
G�����˗�����2f��������ͷ�o��P��PaeFG�K,Q�5u)E$�R�M�F���!:2�
[��}�_6�����3��H�u�kn�L�0�!�$�����iͦ���s*
)d�1�0Y���o@Cz��-��U����6�qfE��	�/|�9��Z�?��P��$�����el�ƍ@���驤S�I���v�������+/>�]��gG3���7�Ͻ����Iyban:��%G0��ȍI9�(Dw�}7�0�g𔣥��<�K���r����x�a����~|�s���#q�:����71k�c���X�b;��Y��x���G�־����tE�/ğ�|c�cP�	�F
)Lx}><�ګ�DR ��VQG�AIE=F' +!�L�"U�ࠐx��&�IQ�G���t�@&��N?H/n)?�>�*g�b������߀]x�������2覅D2�x4
��rZ�����J#a�l�����`�97M�r�e��@hT=<����˙7�����n`&e~�A[ǒ�J�%�%Ǡ�&*��R�	������
�=]N��}l@����!>&������8�1,f�OIq��$[f�W^v���e�3�b�6��ǿ T?l�ˠ��Pu&9i� l�u*l��@�eh����S����qM�p�;!5�&+|��I4��{ B��D�ÿ�8$@���`� )�v2� X��;r�����2��|Os]��A�Ⴠ�M�$p�nw�\ÉPЏ93g�8���W_�@I�F�A���#@���^�w�������ڣ�8�S���0��V`��g�!�b��;;��e�}1 �`�D�gW��cfbnirb/�{[ �#M��J��K�+{w�W�����z!Mĺ�V2w]�Mx5��"G]],>��Z{0�R�5������8�!N�0>��z/������Hy�L�J|x�7��l� �;��sѕ�� lAc**�(Q]$�--�ÎF�d�gh�hz@�\K&Q$�,h��3�Qh�:�OEϸ�O��e�$,�-���ş�JC
[��6�$�'����bN��p �C.>�e�����w	m1ݙV��=Y磟��i�3^H|��W+�q%!�0�4'b�W�b��u@���޻\z*�%�'ǥ����=��Z�޺���B�H$�hkG&�B.��	�O�b�EpL��f!��Q(�̠�����W?��O������<��Q%RI<���9���z�!��P7�hG4���W`ݺux��p��w�V�ܯbQ"�	H/�ܴ����c�?���~���p24�Ċ���dMŞ�N�%S�TO�O�5R��������?X�,Q�L˥���B6��2Ӭv��߉286�����(�c��M9Y�
<q�"��	|�3��?t(o�co�3����D�T����d;��F&�Ec�t�h>f̨�-Z�t>��IN[("���֝P=S�A��,2�ib��tޑ%�c���	��fѸ�y�!RV�T&˖��P��TFGG�Ǳ������fDJ��5��w��h�^��?�@����z�?�Į�h�ي�#A'��Z�;�9�a�4��6��lL�"�Y���{���&�������\�k
b�<�x; �ּ���iCa�qPL>)���}�0M���>�x2u�������� �&#��2<٤�MZ�DS���0o�,��x��W9���f	���W� $;�3W,����*���W`���n�e��h޹�If���A4���bk{�u�2�/��� 96���W��5�0��1ڻ�$ �K�q�Y�����Վ�q;��`o�:h��t���L������ *$	��y���O�{���.(�r���HH�u�#�e�1L� @@��T̓��(��x���-�C}(���-Jذa/Z�੧Wadx�c�6G��$�Lk!j90�1.�"ըhh���(�^4řS�O�+r���]]��wa�P��ī�m�(�E.�����A֐eJ�(���h�|�O���A6�8qA��FH���(�~C�s��F����q���m�i*���5���HMuӱ��Wa�nѢ��i*���ԯy`e���O��<��DC]%��^��k�Cb�����z�M'��2����6���܍׳Y"���Gee%;V���KDH�A?#���~�\r������������	���e�*�|�͸��+�u�_s���~-�o�{�� �w>�9�lNA'�P�2㩧���]{�U5�l����TB�4`wkV��"S�tG��D�s���S�(����H����'��֗&?�HMŻNx+ߩ��\�y�92QP\@�  [��n��J|�c�筴�iu2�[;���o��n�ػ��sf�ĩ'���tpi�)�
��P.Y;�e�����VI�b��{9�/���۔�0�� Q�$-��G,�(�Oh���"OSG���K/cמVT��A�P��t3a���݋U�>ǚ2q%�9Ee5�H 7p��x%Ze-t��UxF�������u��<��8��N�fni��x~R� "/�&�^z���m��=N
���M�t
��__Hjϻ[���AMI~{
�Ê��gF��]����r��l��bxj�P�d�$����X4o.J��x}�Z� �9�A���j̬��Q�u�QS5�{��ګ�
L]<��E����;+@6��bC�T΂��mmh�O�7j�ͽ��H
��º"|��#1�(;�#ݻ�m.F�[WTU����0d��V���jP� ����v7c�����MI���$a�:ʊ��B�!�#ʈ�g���Q��� $�Y��S��0����O��J�a;<vV���ά��c�Ј3����ȳ�'��4J�*�j$SL�'����Az
�[�lsV��x�u!Vj�J�����h����o�w;����`h%\��ON��c3��5+�͕T7�\����X� k�Ͽ��b&p�	G���^��AY�������C��R�� �	'T �0,D'���r4��b�+�����ˣh����"&ko#��u���W0�:j�@���9C�#|n���{?t=�&��o#enP��b�����{���v�ZDJK����������A�C�U�`���8��p��b"�`w���2��7��-�t�I��������s�w�W�����1�?�K.��^|	R�O
T��U�/�Vb�a�9�d����X��ۀ����������;�x"�I�{�@ �.M3�2Ǔ"�4�A�l�j���� �M���L�ZҌ��-.�=�(0 Q�,<V�|�#��5�����=��!�J�k'$Ň����u0���SOb�?erE��e49��g�*Hv;�7!�1�dTp3��*w�D�;�� 	���D�E��x9t[D<�#3�#�9:oF�Q<��l߶���h������3;��A2mB�"���6	t�0l�����&(L����N�bJ�/�E��bFS�#e����i]�6�ߔ(�P�� �]�� y� ��$ r`����9$�)]ӓy R��m��w�$�>��#��" 2���4�Z���KZ3��nyެ����b���N�@�>7�p5�5X�!�Ҕ���>�z��� �>�zjO�+�u�^'�L���-���%�}0�W6�b�hCi�S��N`q}	N^X�e�
��>v4C�m:+
ʦ��1�~����to�O��E���h���(@�8��@+��GQ�
>xJ��+��^9���I8���PҀH��-���Aa`D)�	���j&q���K�Ĭ� PVG�[ ��[�g��8�u����ס��@�l����G8��Q̪��џ}�d�%����k���U3�C�N�c�@���%R	��	,��Fֵ5�P�~�(���(�Q\r�r�qӇ`g2�Y�����|���s|�
*l��Sה�c��D�����P[Y�.X@�T.�EA${�:�$�3NX���z#4M/���={� P�u�GF��f5��H8��#�i�64/��[��SO��;BEa\�8�����&zϝ�Hعm��������BOw�344�eG}@x���o��m466��+��+���g�y3g�b�ѵ�T�w.���,��Ɵ��K�ʕ�\z؂#�+cdyڔ6t�߰��
��~+�53�?�D�$�a�]��ʥb���n��9l�J�"<4P Y7р����C�"�'@41����i|��C,z���6�@o�`�z0�hI��C��L̘1G-����r��2 �s���B�g�SD$c�< �cör�F�VaRē�|���p'J�ȟ��k���u���H�݄G����j��`��������o0󶔖�񄊞H:��w��dOk'�E���=A�1��(X��R僷�&��P'	�l�O�i����P���زc+@�G[��P�a>�#_�(W���Uo�`&ym��\�
~~��ӫ�6wr,{��:�(ЮMN&�,�F�urp:B�n��!��aS9�E���8 �2�T?��R4oقl"�� �:y �����S�����߫SO�Z��[���g꼘Z�I+@9 #1�D͏q�B�@}��Cq��MN��,�Tp��Zՠ�D��]�#D�Y=QPPR;�]x5D��]�Β�{[�B��s�k�i��$��ItJT���0Y����7`�.ů^�D���Q$�E�D���'\�Np��
?O.1�5����\r�)B{߀3��Jh;0�̚^&tƜ�J7�e`ء"�)��zg�s�7~�����i��#�M#P`��hz1~���rv����Mm���DF,��&�
T3M�/G����QL= ���	�,3�F2������˟�����x�=�|���1�K0$k@L�Հ��[,��AL�UU���o��2�����Ғ��Qf6	Y���z����/v����8��0��{z{��������A&�D����Y�T�я~�Z*��>�<�z�H&R�HT.�sϮ����㢋.�����
��ҋؼ�M~q�8p� kP��O�#g"�5�t�R\p�yL�b`����<UVQVaѺl�A4'i>���PTQ���G�R�,ƾ���!����I�Dy�7G�Gʋ�s�����=�?�����":#�r��?4�Da���>=����.s�w�uz��A�&�H��'��5�	3��8՞�Μ� �-�m3�H�c��FNO��C�FR��	�x�c;�$�n	~��X�LE5�ʆ٨�>��4����&�� ���IS2M�|� �M�c@�ɦ�h�"��� K`<��(A"c��Cz���cᅑs ����V4�5 $>G��WQ_��/�%Z �?�d�,h,��[���4w΀dq���!R������@) ������Q���t�+Zd��L�~��ǘ�) �(8����T���`�s
�H؆�?��a�ey �q)�4�*�4��̟i�U�,)��歈O$Q���|��ES�36��O8�]��O}9O��{y�.���ѝڷ��
�tp���aeM莈����oϿ��Y�PF�d�@N\X����8�o{��`�\�`eN�������u���� ă,vn�+�;[�d����T&M�B�U��"�r"���V�_<�	���8
Y�`��2��,M��8��Ȳ���@��2>s�Gq��up�vw�9���£}hșYqx�}O�s��7HX��+`	"�~	NfG4F����l<���A���Η��F2*�9r���w�:��-CAba�
�{d9Hy������7^
+������@���g�Do�A$H�i��!f���S)���z���9��D��-�Y�`d�X(	�8����g���ak����Ń �?%���bEEٙg����������:�8�ðL����H�3�e�er�Z����=�4&�$�e.�J$Sn�4�>�y�2���y�D�;��0w�\�K�|غ}~����Q
�,R�"���3��4�:�`Ix�Q����󖢽�pH2�{13	z�T���D� �R����8��g�JT��\~Y��ņ>)��>�a|����[6os�GF1<<�:��{���dQ.f
ִ�J4M�E��yNS�6�zz}
�/zt EQ��F�/���&ED��BզpE����>E��H�t���!\9�u�Hr�K�$X����Q�Z��ƣ()+EYE*��xB`˗/�$���.L$R�V�td� 5=k�
�~:��6m��Y��L"��iU���K�$�x�����(2��Q��)�s� ����
dew(��x�끄�v�~��S�
��P�8<��n��t�*��|fo�$g�´�0�	MX&�}��ȡk�m�Eع ��e�H�9�5�<�ȡϣ�i�ը*+��-�lGMA�t��~ӵh�Pa'Fp�1S"�������V ��ja4��S+�m�z���Q���@W|��֋'�l@_�F
(g G_�^�/��3��el7�;Q$��{D�S:�e�8媏B�.|׮���VGSXB�����}%��q���C��@W� �F�J#�#����Rdߤ�E!U�%M�ɪA��ܱ���ëIP�s(d�h�ꊋV�����a�R�0w�l�r�����N����Jؓu��z�Y�" ���T;������wɱ��0��&q�7�G���x��#
d
�ˤ@9J��C&,6���9X�G�vj��_��G!�&��e���O|��HIE@���]S��������B�-�FB�Q;���$�6!�)E�
��priT�zq��Y��K7bn]Xx�駝ʪRZG�h�+UR�����ǭ@6�����)�䠫k;Wh �	%pSQF�^Ե�U	�X��4�4e3�2N���3���(9��й�&c:V�f�DMU5�*�1g�\87lF{k+��T�UbfcOI�j��[�����k�cͫ����}Ř޴�4�Qa��P �#9|�}O'Qr�,*9�ڡ|
7{����(�!
s�G)��L��sN�G�� O�F��X��������Q��N���s_b�$�[L�>G/]���j�}L�F�L$��{��j����P_D��1%�։�H�M�F��Ci:4:Wl��~]�A���    IDAT��� j���jL$2H�s�Ch���c���U�PU[�#/E���p�^��z��x䗏�ǝ�s/�O<�
�75Cъ`t��˒e�
ez-
k�ȤiH� {e��{��)��(�C%r��P�H>̯I(W���x���H��<���\x'r�;�}jҝ�o�{\�~�=��0B@g 9h�$�5�$� Fh�A���0���Br`�D�����JTFJ����(4YF�&�֛��5 vl�p�vo����9��S+�]�����bS�O�@gw�C�4�����9 [;���s��5�4�s9�jV�+���ዷ�jCȓ��8��8�ʫ��TC�ߕkm�o��*6�n��?�$SGyQٌJ0�x���ގ^��0�2
��s0M�mCYs�:�I B�j���;�"��,�B�B��+�"��
Z���T��!rD�9���p�gaV�,�v(�cN�/<�k���G?I}D�:rv���[��	G�U��ux��?C+i�H�r	�P}�\�z$�:�ߠ�-*(���e�xDh2�Y��Ÿ��!䨀��ڇk?w2j1r�K�b���1m�2�TTD¨-��kk������f ��+d�$e�(b̪�Dcu�q��1Կ��ƀ���~d�L�ص�m,Ğ5k͟�f/d3Lɢ4������ʿp1M��Lh�X��I]Gq�7s)$����$c1��}��+�T�OnHE�!^Ǫ�JTVVpqM����$)�UUT���N´�:��ͯ��46��W��M[��Kkay�h��]���`��|�DBiC.ŅB�HL�Q����G�Ppp����BD�t2 W.G�c�R�hC�����أ��ٍ(�i���� �;��H�000���^����u`<�cPS]��"��^�_8c�v#pES��ߋ���B�$��Ni����E����e�Ih����8PU/�XGi��M��x��C��"���dI�r���BO_7j��0k�<TU֢��������x���q�O������'��_y{Z�AU&i�|�	���i���x��L*/��ȕP����@�%#���U�D�z��h<�riSȹ��O6\{ 7�q��o��y 3Y~�[U!�$�&�MG��
*��������6	
����G!�=Fh�	�s�"�)P>Q�
�7H�S�{- u�غe��1x	��D���kP_*Î�SN|W����/٩��Z��
L]<S���
LZ�֮n�ɦ�pd�s@�u�WO���#Y��LÂHQ3�%��8�3��BKw�HJCur��L��.�Zi%�лF86�ˑ%�c���o���d"K�H8R ;�t�,�,0�Re4N ���EX�íh�O�\XQ��T�����L��gRq���E���"�0�:�9���	����`��q�-���ڰ�w"��-���|��ǎ�l�=�����w!I�����=�g��7Fi�BLdL.���s�g��]�-��*4�!���}�**S�h�)�M������/FC^�Bk̹��wbD���hLCs��K���$VYDUI1�j���aRB������R�MX�4��cn}%�4Ubnc52�	��,>���m���ݻ� :�c(	:�,������Վ;p���� ����l�,(R
����AP�œzMmu�����)��
����1w�L��T����4��Fa��7l������QVR��>�e�8:�M!�g���s/�ú-۱mGԢr�7�E�Vx� 25�`�u�
��Q�J"n1��'%��~%�z�(Y��Jz�!@l@�P�a
G/��Yue(@�+a��9�_6l@*����(S�Ȇ��W�Cî�%�����A���p�Aٲ���k����v��1��J6��l�IG#�{�h�HXnsX��	������ƛ۶!.�A
v��lNa}д04؏��.����c��<��?o!f̚�D<�u6bWK;�}j<��X�~�Ƒ�ZH$t���Nl&	��^ȵ5�%ry�2�� �u^��א�k8Ȕ|�2 ����Y����țl���W+�=�Y�
@�߬�d{[ ,����a#��y����^dkN'	ӂX�DZ�$�Aă"r�.�Y�P�@�`��d�Ţ{C�	�R�D���V[���R�hފD,�"��g��
ӊE��A\|�IS5�T1���
L]<���M�콹�v�8�LF�@�v�S���3�߭\���l	gcx��FSM�,��QU*�X<z?��	*����;��*H�b��w�z�����d�x��_  �&���XNB�Q��杈�"�`�hڋ�x,�_�	���p�0�}O��, �N59CQ�J3�W�B�D����\��&M?,�>J"'�7��@Q���/8�_|��
��9�� ��ל{�+��a�jL/��w��dŋ��n�=?�%t�Ѭ��*�� ��[����&-l���d�-�e��l��t\q�����@�̈(��aǹ��;��������]\�-t8��t�P_]�����d�G�I�(�]���\�BڠuX<���cɂ�*T��� ��I�\��u� ��@yz����\�S�H��T7E��Y����L32 ������v\*ѭ��C�0�iO����"�I��p�
�U�����x镗����m�i�eU8r�b����XlM��a��W�y�n��R�M�3�H���I��il����g�h�4{���!M:\j�7  � t<�k�#:'���a�N��(N=���6��1d�E�DG۽w�*k�����>}:�lߎ��>6��`?��Y�Î_�H�d�L�V���V���rZ9�f��SYx�'�ؖ���O��	�i�A�G��k_GIi����d�t\	�h����Q�EGy;��D��E�^T���_��}C��K�����ֶNwraQ�9MB��\Q	��Y�z"O�h��g���"z\Z^I	��4G�od��Ӈ��C���36� (h8�Pg����C�s� @X~��žه@�[�BX �h~Ѧ�A�ݢ���̕�������N _����:�
�@�.<����W�'>��FtN�!�)�j���E $O�/yPQ�ŧ���%��0.8q��Y	L�տb���_��S�1���
�����u'g!mH�2�F�x��m��;C+�nؠ��Gi 8vA-���3ւ�7���Ɠ/t��^�+ ]��ozG��tt�#��Q�F��¦�Et���"�tx<[-B<���뛑�4��2��$�`o{���)0��ҧ��
)J��$dQ�iSQ.B%�{&	;�G��84����
�h�mq7�����PR�Hp��Ee�u~��;_�*�ȥ0E���Ꮋ����b��(j�^<��C���T���p�goCF)�h"G�pa��Kv�n���	H%F!8&gv��BTCn^���>v�i��Cg@�Ǹ��T\{�װ�w���5���R>
�(V*�#��� µ��`d�~X�4|!?�9��{���g�h��Ŵ�0�c}��P����nx$���QRa*�afP^^�e���*u�ɱ��FN7���9(*�*���N�r������r^��1�t�qb�$1�!F8b;�L:Ɂ�A����e�Q�\�0%��H�2x�x䢥L��lG��}�9RY#�$&�Y��'��1o�Rl۴�����<�(�I0U�)X���P����Q�<M\���9n�I0���H�ܳNƜٍ���_E�W�mdxb���#PW7�����Bq$�Mo6���!����S�\���T�/�[f�`g+M�b<:Yrm�I�Ok%�2_���4�=�f�Bǿ Y{#������,)�H��wo�i�u���`t�9.��BO)��{ �*�x�����m�a�l�;D���녷�:M 
7H:��7-�>U���@Th�x���a�2_����0Šܖ�$��`�+J��I.VxK�������R��˻R�?�8�ۖ����:6�L�c��.��]���,���i^�}��4�%8�A�D��$d�iȪ
3����"O/�suʡ�lv�#�ʊ2�UT�=�@� �?n��r4�)@z�7��n}O��{ޑb轿LS{����;�,g��̊��F����عoN��s@T�03Q�N`z�@�G�*Bf�u^*�m��B�4��Q2c!�;c�nql#��� ��}�ۼ={PT�LƑ%W]	Ƴ�Z����E�p|��2l�v �Z��n;�x��N��d�I���Hk;��>��
F
/�~UA����۝�.�
�U�!yC�� �uӡ��P%>Ճ��~�u������aQH�b)ǔ�x�O/�G�<Ơ����W����"l�p|������yz�uȡ�4u�ɹG��AQ���bɂY8�Y8���a�4#�)�]�ʦ٬I���K��/�f���귯�rn��w�R���^.��.)ij$�)�BA �Ē��(x�ٕ0ƣh[���E'�&�����y��Jb�ڗ`��H��<�pu2��#}>����رk;�Ϋ�j0mZ-n��v�شr ��O�%���|� M�20$� )fc}������R)�Y�U��8н���a������� ����4��U�#O��"���Qr)�Rb�f����(��Q�����<A��Id���S���'� �F=u�EM��Z��
P�-l ���tB�b�;��^	��(J��8/B������ K"�G�9P�������9Ẫ�ٜ���9�o� Y�I��Y�s������]����琈���Ņ1[睗L�*Y��c�w�4J��{<,�&���}8b�b>n�-�����+����Ǳ$A�����������0T_�a�5M�DÖ�j˂��Z���_ ޲r�ug��2��LfJ��HZIfڢ�b�v�^��f���<�����E��5�1���O$��F�����$%��ڣ[��賉FGZ"�d.���sYU���z5�9�u��#�'��{�ҡ���D/#�92} 3N}'#ivx�s��H��D����@Mi)��܂T,	UpP]����r�(W��M��c�����]����|�W`��yǗt��/�@�νN"��"W#ۺ����?1X]'�K��M�֓(�28��\q�2��4s�J�,d39�Y��.������57޷�Q$���\t�;6a���(-
���8y9aJ��X��]	���H$_��~ )�_���˹��n�i�<jI��G������lY��Ň����M��'WÔP#�g��@<��F���?�:�6�M�1?�Z3�s����=�XX���b��F<��]�����T�����}��[��4_��� �X�.��K���7��E��H$- �;�b�T׳���ⴣ��7_�J�!�~��6�s_�6��M��6�����;�7�*�H'�b�2x�{�n�Y�	�Uu*�xs�V�(	E� !'<6 0��c3���fpd��8���Yv���6AB�2
�N���Io�|�\����׹���#q�=�}�	UU����{�a�˟�����e��S .��n��ݻ�#h�`y�䇔���T�G{�����*>�{��Ǐ�Ѫcrbc�*������e���	���8�~��|*��J4ELh2�!t8��-j2��a�+���v�NK#��b��3�
�|��і4�H�bN�P6SJ2�c�:RÏ��'�0;�>�eS���hv}Dlś��'�^�S ��E/�ZD����L������M�ê3O�b �ʝ�.E�����}�RAkiEϑs�1$���������9��8{���ϡJ=K�-���n�+Sד$�*���;�����L�W��98Q� )�bE�Qi��$A���wɶT�#b��n60�pY�+�ˮ>-��F�M��b5�$Bsc�n��H�.��v��H�u�F�d!i���1�MϤj�8m�,���Ʀ)�b�L�aU:��Rx��72Y���K������8K"�����h� �@�b29�܎R�"�?ך;N0h���אN9�*ze1^�v{>|�|z��`��֍�`��$�=�'�a^2Y�/���c�+h��/��_�}�L�_�}���^<�����Y�{Κݞhni]�����?������L�p�Eg�D��{��_}��t�^��E�I�,�l�C�ӂSŶ�\���� ���M_wq�X�n�b�V���gO>�եE��R��"�@dyXh�x��"άD����4V{&�1N�Yk-�rU��"�~�,���/;���nH���Cw݊�֛�Sg�3R����0~�>������3�چ-��� �#r�+�/z���
[m�x��B655�|����<)���s�p�)|����!ݦ+�vb�?�%|����b�� Ķ�
Z@���W^���?#%�u�j�������v$v	����ꆫ�;��g�=l+�hg�g��x�a#�]��:t\�AB�a��m���dp��q�:���%H�z�o( �nY�n!`D(��4��3�3��VW���{m�{ɟ`�{�34 ǲ�X*���uUV��T�ҥ�D���.�1��5=a�4�0��9N`h�+�g�)�~��W�{M�� eo�}bw_��,�	\�H���=q�"�O���`w��FG�S>GS����w���$��t6H?y[�8z�!f�{��B�B<@5
�M�	���k�R++�'`��m܈M����������p�h��)K����E+�d�?�c�-��Ϧ.B4�rM�)Y0H�/����jt���d��+ؼq=}�Au�$�� ���$#Hpq9Ւ��$&�ZD�@j��dd�:�h�,�pJ�cc�Ŋ ��q��x����6�sGQ�i
��yǉL��)���
����;��G�ڦݲr-����4<�$e����7;�A��˨�\��_�4"�d����J����bt�=�߰����ae�.����tk6ZB�:��*��+��18^��L����4VWV�UGp��$6�Lc�C_C�Q���q��w��[�k���"^s��<늀�}�V��.��m[8���
|W`��G�F� R(��������;��P���pӠC)#I'��_<���~N�*i5�'�c�d�H�2�25��^�J*@���ƭy���&]���,�Q}_�����"8��N��6��8�\Ƒ3�6�i�^��V�}���jY��W(J<���(H���I���!8�y��s��G~x~�W?�}���1y�f��W�\�ǍϿ?����%�S�t�kϲ�K�=�w��#��E�i���s��DOX�.�3
�����q7<q�����n�h�m��n|��x����w��Ѷut��%x��߆��,V��i�?�R���~�8Q�e[G���w���>qq��*�8��x���^Q:�<滶n��S���c��`��c�XG�+I�]��8�C��� ��F�1e��B�*S��n�C�т��a�N}q�����$2Ѱ9���B�A�����X�^�H����	�ԝjv�#:�� ;�|��G�!VG��~K�*�X�܄#M�)	�^h^A�<��S	<�@�x�\�k #/�s "�{1WS��9,N�� P�B�"�K�	�R�s\Ew-|�JϘTFk�Kb�@�^Ƕ�۰k�V<x��X!u�6�a$V��uj"41[;�iP$�|��M@�m��Ш׉GA����5�&,x#�(�F$_�z)�@.߽�~��%�ᄮ�U����''��"Q�I8�EԤ��1���uQ]�~� E��J��.�;V��
�(�Oq%�U�_<g$�&�;1w�ʏ���_���?�z1���XW��\?N�x�#x��SV��_{��c/��]"���RU��m4Z)���=��#���`h60���n�j���'�ca���������aF�����;�l�Ʃq�}���uQ���𮟻;�*ڨ>I    IDAT�x�K�A������e+0 ϲ:ܝ�
�}�HVow�cL��Nbbϱy|��#8xjaf#�]�]SR!Lv���x��\�]3԰
'j��-b (=F�ư�.���zG�Ppk(M�'���U�ìw<3�jD��a*p�`��@����N�<��O��`��Q��*b���8>��.�M���Ml�Ҫ��?�\�OW->�X��.v!� t�"���'�����1���Z���й��q*�6Y6>��G3���	]�z�".��k��f<�БRtr���<�O��q�}G��3�&'�$=D�%��ï��n���\������m�h�H�����f#�\[I:��^LEEr�E,�R|�o�_|��Q�N�q��Zu�p���G*���ܹl���_��T�q`!�m�5�ٱv�m�0�L=>}�C�[~���6
��x|R�:�(@ub�nC	�Y��D��m�e�ᎎ �LI7�;7o�	ʓ�/"���g�v[�<t�E��a�Q�� ��24����.y�g4`�uPn���q�>t�)�*e�ū�!E�B{]�fn��� Y��{1�CU��S��\ù�k^���Hz��Y��U�#�p�^~.`'U��������)�6�wB������X�A;�lŎM����}A������ D�i��͂�B+YU��m! �k����M�
����O�9�<���ĤLc8�H���v��o�W��_�clbW\v9y�Q�fr}R�&�B'���VIaQ�k(J.j���rtR�#w�˧�8\#`�xh�[�Ra�z�#4:�)�*������sU~�t^�L]�v��Lt��v��PV�l�t���,����&j<�)�������W�2��RĨ�)U���V��N��.�Ɠ�,�U2��ϴ�������c�����M�N�PՍ맱qr�D�l����W~���>UBԘ��_6Ԁ����W7���|7���
<���l��Qb�r�����W���S�R�@�E � F�a�4��:����c�r���%0�Bq�9I 7?3)FH(�jBu�ݢK7;�A჉�t,j�,���Q_�޹�Xpl����p�q�Q���K8tz	�	bg�����r+��J+�]��KX$TD*��p���(ǨL�`|b�ɮ��N�<6�Ruˏ}?^{����j�T	��n�N:_���J�z�TU�k�[�?�����%�R#�;�҉�TJ{�WH��q���������G���c�i&N�t�O�p]���*����C�z������	gW:H����4�$�����1v���m��ujF>�h���b�E��cƓ˭��һ�k����~����ŵ;w�kJo̺��t�2e�Q,�E�Az��p���G������Řرa� ��̐x�5נ���}=$�v�*��l��T�ґg~�G5�$h��̇5*A�y���If�z�ܖT&�θ�&t��t)xj
�_��$���ҮhU�&R��{(�[�*�sw)u��L��J�B��#r��PMg"���SSw4�Ie�%�E��/P��`�r��<�m(Q�x=B���M�m�&���O�1Mqc+�K2Q�6R0���ETl�Lb��p;�M�H��i���b؝%�R�F'��R�g�k����=�n��.�Ka$�h�?���=�!��IJxB�0bE�c�A
e�u�3*;-��M@���_��R�Kޏv��>��H�e5�T4��𿋧 yN����m������y!$�"�N�D�715Z����F��7���&S�$�(��Il ��>jiu�mI���� <��f��J�	?�R��:|m�g������p��"��ʣ��\�3��z�z<v� :m_��S5���7a�ti{	�{��5԰���7�Ë�\��˞�+��Б���RdЫ�c��y�y����.U�ٗp.Gĥ��,>&� �֕p��l������UuM���B�D�s*n2屚��������9�RC�o���gq�l�Jw�7i�\����@/2�M-<z�4�}+��F�"0+h�zQ�mt�̢�E��69}�e�!�8�~+�xy��K6oA7���H�}�p��߄�ز~ox���7�,�#��q&�5F�$U!G��U@����3����­_�OD���,�U�$��p�L�nv�¥��/��y���q�z�D��1gd�؄q����Q�V7A�<�+�<�Cw{��/~KMG�. skH��w��mX�:>��^��t�wߑ�/��K+����v�m�������R+�=����z�]z�KE�R�B�DKw1�@���2�@R�)p�f���Į��1��]�$�՗]���
�!�,���N��qt�m�b��>Je���{��9}�s�U�[�LH�ʩVR��tD0�QDԲW
 �D�㤌���;2��y���Y�����8�����E�"�ʋ�<�Ze�(q�������`B��^����鹀c���S&��G�na��M�b�.|��Q�# ��f��yK{W;�y��T�c��K��fx,y�ĜB�Q���	�PT6����<�F�Q�V������k�ė�x+�vO�VхN}�2�p� D�u|B6��Q�C�����6�3�J3Bj���L��DVUk���
��M7.�eL>�W�T;Y��KE�=OJ��౼����C��P�%��XY�]-�����u��L3��z]a�I�#_��	y}�Z#^��$������=ܰ}Z]��,k����G�����W���Ԃ�fB�H����q<� ]@���!tz��L0Qqe�kҁ�Y�k^2��<;+��^};V`@��<��g�
>y&[�7��Sݬ�}'p�#GŎ�|aZyR0�b(It�Ŕk3F�[�Ʃ��|=��[�A�Ҫy�H���|��Fd�4R��5�����)IŖ��f!�~$4�H���*sX�Ć��N�'O/���V�E	�;�f�!0�8��D���ۋ��%��x���
���l::��Fmzcӓ�Em�=�Bq�%�B6���o�hǘq�=7^���x~�y���'���^�u]�ߟz�x��?�o�[ic�OP���W��B0\ؕ""
�� N�C�\�wP�"����
�}�[�e�u�	EM���������HLO2=��XmE�"T.WЭ�`�b�{_�B��G^���t[J��.*�۩�����0Z���72��0�S,`W�0�>>��~�W�_�CpFfD�nl���'K%�t�e2���ra���m;��V���=��+Ыױ��{f��I"3چ��c����(<�K����8*݂8a�0�Z�~�J�jx�?��\�i�{n�I��d.�"��IM�8�P�U���^kAp�:W���~�i5B�}�𽤈�* ���X�k�:�@�RE�g:x
cl�hVف����˸dz�7l��w��ݒ�k��ӄ�9�͊�'�v*N�]�hm�:��&�+чm���u&��&5L%z�ՊP�l��V����q\~�n�u��@� D@�<�͔�!�!����(��J��3;�9�orR��ܐ��~�x��9EJ�x\���pu��<�O:���t_�}�U���4`R�<e鴦��
��j�E��ϟE��0>R��m�U�K	��v����	���z6Ο?�2CG�$߷��J�evz7��Ex�[��Qa��fׯ����}����Hݪ4�x�mڸ�&�p��A4ڜ^����?��[�u�@Ҙ����E��swn�w�
/��#2ܞ�  Y\i�<H��Pā�K��=p�\A�bFY�������2	ϸ�`�%#�b�86���jN��`���(�Lt&5Ñ�Gn�1]�T����d��U1쪒�I�ݴm��F�[n�șE��"����A�a�k���D�)i��m�9dӄbé8�R�1�L�#�-�--�p/�����i���_���D����/~��"e����OIE�<"��{�}w�y2����$-?��&)�J���6<��H�����43�7���a�$�$A��JFϝ_���U��ů����Z�bm-?A��)S��A�5$AW^�֍S& �j�Uh��n8C�O����$��֕]�b����u���������`���:KK�P��6NBH��Irs� 	]O&jT���碻��=wߥ���!$-��Ӗ C5����"nD&2����J	�rU�j(x�gu9��hJ��K��[;>� ��=��R��BZ4"�>J���}��ϣ��NQ}�j�A�@�A ����dI�AA�`ݟOFr=�.�N*"-n��I8�5��2:QO�F�4D�n�bZuK8}��7i�03d���l�Z%sG�K����?e{rq�^����E��tV�%2��Ie�T�W�`˦�8��C2������$3H�������c�@�=�x��$���W��E��đL��kx! 1�<�Q���<E���:�d�<�d��@�4q�◛8~100�]&�$��u�i�Ŏ�����`r���S2�#T�%9�=����͏�j�|��%8բ�Kw��O��7⺫/A�`d����¯��`��`y	>�U�u�&�߿����~����;ފ�U X>��ŋ�5Կ�{����^<��7����{�x�������{`1�pw��o!Jm����Q�C6�̰b�ڊ���2$�<]�uۦ1e�(�jv������lF۫�ha�QP�DB8ـ����:AIf�XA��2�(�k���b�����nl�P�E;�ъ\�FK�N;#�J�)�X�]��s��0Cu�z�l܈F��F���t*�r҆� ����t�2Mq�J������ژ��kY&4w���HΞ���F��8���W�&V:���Uf\��+EO:���E�����=��c$R��~�JUYj6��L���F��b�bU�j#��@ҽ,��E��b	�r���5
��E^�7o®�;p��	��A�n��q�)����X�r���,hI�b[����aa�K��2(�R\w��Z-<z��LD�TT� �++�\h. "`G܊Xl%���\�A �/hB
0�Ԣ5�S�3Z�
���Ҹ��ͅ�m�r�2輦5%kE����)�  Q�rNGh�p�ܧ����bj�� Z�-KC�F��`�9���q���A�P43I�O{>� AX��z�_@'�}�1' g'�s�|���(�.�RY��}KK�,��ѮWk&�k��<����85e�����_ydD�P�Q�qK��&,���U�ȐjE���s�������q$9-~�g�@4y�� 5���8D�-���|�i����285S:���581�_��:��� I��+3X�Qb�\6)�K�N�����X�&Gg�pr�g��X):��B)Һ:	ෛx��/ǻ�'q�B�_:����ۿ���=�W �ƍ�v{���XYm�N�����o��R�����UC �o~��w�
�w͡��7���9�-7�(yl���	��8�/�9�'���c�s4<e�73a��)�X($� V����"�V�ucULUM�X��Jf(��������95�H���G��H2S
�6��D/1��E���\�k5���t���L���U�[��x�V�	Nc�W"L���a� �c��D�DR�hcI޿PA�s�r�,��dij;���К]B�"�Ѫ
�c`�d��ܷL�]�.I�ϔc��+�n�*�;T�Y���1���g�P@��4W�AHk�D
u����Q��2�ˆS)���qO��b�E��>j�U�I��H;]�� Q�y�;\�UA�_N J̚0-���Bբ�����{ �yJ�
�<�L8�IL����;��͔q�taǦ�(Z��s�tݹ��r���*̔�_u�9��TF�O}��	>�����ȶJ+�s��������H�*,p-TO�����5Q.K�;C�3��`�n��Ŝ��ke���,`ȗO�����+���DE��`��	9�i���e��:�X��=�XZq�2S)�,+�8F�䉠���e�f�9w!5<�
F''%��NI�C�%mO+SwʔD�'yq�uO8��"�fE@���	���~H������94��*��-� P�.	.��K4IZ+#�-5����Y�@�,5up`��^/�~��Ϗ�����5=��4LkF���i�\羑5T.o���$�NQ��H�&�;tG����^(v��W��Z�Ɗd��ނ��hb����'��x����G)�l�& ��G�`i~�r	�'����}&�Y{	?p�M�����3\��Y���3<-�+0��;�-��-�WB+���᳸��8xr��H8_�z��قe(�(��>����g�e��m��������5`܋`�0�U��	����K�,�e�n2SR0l/@��D�j' �KD�(��F�K�^��ba�)�v�u�
�NF�b�%�@Tt�=�6n���Z���"��(V����́\3�2g����yE$>-�c��%릦�
W���u3mC��A�5Y,ʔ�����*q�#��,���Lۀme"&旖m�JxM%�N���r�I�(�����R��b�B��"�1.��Z���N�� E�$f���s���(OM��"���@���<:_�Wj���૟�<Хm���e�������L�؎�U@�A	b\�c'�vzPi �^�,�����Ob���A{عs��v�qD�.Jcc�� �/ ��� ǒ��!���q�A[�V��I
S�z����P4 �g���f��m� �j��G��X$!x��Ծ��>w�9�T �lعn��3������e$�) .�n数�g�;s�u��ފ��G>x�3���S97
6;�*�$��T�,�O:�r��܁@{�n��mԉ(`��qE1��bZ+����a%ߏ'A���(Xj:+�.%.ρ_B�� ��ə'fkz�\��O���n � �?5��\��ϣ�ϧ�\�= ���`YL��p���,�m��/z� �0
U�G�ጊjh�6�N׾�ض�|�>#�W~O���ޯ�/��z���c���}�s(���u�-X?3��{�`eqe���x���[�����:^��aȰ���7�C �ͮ��u�����q 䁛�?-����q�gq�%���})�u��S�SX�*
DP�[������BeԊ&���b�D��G!j���5B��T%B!a[|5���J�Tfy���ًd�Ed�#1K�u#,.�1w~I������ Ee�ʢ,-�6�������e&� A�K���!x3�]��A*�1�>	BD�H)삇�ӕ�S�E@/e��S��#Մ֒��/1פ"�dg�f( DuJ�\�'�稘����B.Xl�0YhH���<-�S�n-�}A-54�zkN#��O��i��x�z]�+#�:Hۤ���OS�4B��.9)/QbH�\ɱQH���8�	�����5sm�N-��܎�� HRq�}�UWI:��{���8ƦM�q��9Yꂘf��f�ł\�<Z M�#�i4������.$A�yW�@N'�_0��Ms�F⚤�Y%/B��(�'ҫr���$/�s��_\��s��s��	�
nqI0�HL[wWMed:@k��P�Q|_�� ��fb���adrK�:P(zp�B��!l� k7DП'�+W/E[Y+s���F1�ng���l��{��8>��!s,DLx'0t�tω�P^��Y���� ;�,��'"����u.�Zi��׫��*�\����)��r�<	�����=����rҨ�J"k+�{4�ש�t�x�I�Ӂ	ي܊W�M��������� $�Y�s.���l�%�rH�&I��vWS�\��i�V���^���j'���1t�l�����k�5;��˻�s�%Ba}��M43���lݲ#5xt���8 Ύ���?�l�*��x�M��P��J`�Sߎ^<ߎU~�3f�=y2kt��iO( uʸ{�1|�x����1o �&� 	���4֩�,�@�<��4E�=3�`�\@ձđ����3ک�0�6�$@BZy�JZ �	�v��VQ��%V��B    IDAT���8��zK
R%6W7d�����t�aǐ�x��)xc5dBϲ�nw���5�(PQ΂����t�H�J6��PU�*�4���%�j/$�Z;��/Дv� gÒ��ܲ@i#����J���O��%\x���޴ SkFYor��;R�ԧ��TXdb �N5�!�9A#@f��J�|bb�OϡV����p��M�v�T�p�}(=���G���0� ���<�ջ�&D�?p���.��%c;w����B���^��3�qd��>��������O��C�f����Gu�� <�n�n�
uU�����s�|�y�g��Yy�.V	���y����σ���t����n]�}��`d��Ĺ �b���Ą_jd���E��dV�\t��]���)&<�;��������!���N[l����u�m2$
�z�IJ�+�lĩ
��vE�n8E��$ةhLy�x��ՠvй�����o��Η N�Q嚖���u�ʟ9@ �N�K�e)RY��sX�)դ��#O�P	�DG��p�߬���a���4��CMD�^��4���󉙬_��b91T�Fܰ��M�wB���~꣢�	�R�\���wBW8��Qk����Ce�Ga���B��Ƈ����w����Iofv=f��qp���к�*~�m?��3d�U�|�����<��p��^<��R��ݰ�:!atLM����4�?���^�\DgA B�$���La�8&IW��9	�S��sf, X1�����zX7>�j!���a�Ks���N`�bWg���H@�u����A"���|vș�.c�: ����be)�C�ܑ1�˷�Hr�&��쒊p8Qal,�#�̔m*' �X	��!1T��z�SzX|S�/����	6�r���Ԉ�K���@b��s�F���uE�X�Hҷ�ɲw4מ�?�U�XW"V�����&?��x�儘�dKK��۹m;�<q��i�UI�I�^�2��M<vp/LNJ�L�"z�20������w*Z�$c�}�J��8���]B�b��}ΥX�_��GV�K�a|b��Ә���k@���!�A/�u�e��� Aw��l��;�j[�� w<�Ԏ@L��T�
��R"sE%��] @�\���6#��*hj�~.(���S�  $�4ZUb�N��Y��կ������.(ʙh�8y���±�.���� N	�_sݩ�i7�<k���Z�Bܤ �פ�d֖��9�&	ʐ��h��.�JY\��Z�煡 ��L.9����B�}�'zP(�sOgM�R@�ǣT�����Y���k_�a���	����m[������ �5��� ��{�y?H������Q�o���mU��j:>���u�ב�R�� 5'��Lڤ'�#�b�`��
��DՎ��>�Պ(���'�8�~�q��"5�ܱ��2�<�4��C�89����G�s�����W���a��P��[�Ë�[���7}�����?����a���^{����y/�5S~���9A�:�SgJg!7W�ʘ�a�Įi�#`g����e�4H�r:� ���&�6,�%D�!h�u��&蠆��~���B�Z]X^I\r8�����C[�4�U`)K_���F�0�~#�uąD�((QuN�aFI�-�����]DgI�3��pɶ�h�-����EX����5*baKw,�,85��ty����(p�����v��s]eT�tX����-H�n���Nh���8��Y���,yYD�p�Dv���>�\s�D�k�X��׽�5��^����s������Œ7cX^��')֗o܄���u���"�+�?nb|�n4%������؁��
�< �0H��^���(֪��j	�v��(�*�i��&��J2ə?����T42q�R�%��w���ZS���Aҹ �2-��q��g�6@��讵L�X0j͂E���62=�v�%�ϕW^��N�@�]g�V�� �vB�#��Lnل�n]NK�T���U�� z|�������*��	�Gk�@�X�#��|P3�ʆ�9!EO��RG[u�/���h ��m��:�Qhާܼ|ʤ�\
l�`V@��J��̰e��f����Q@#ϑ8^�yp��=_���Ϗ��p¥�ok.Zk�ŅY0�)[.���ާ��e�"�D�rNI��
=mR�r��򪅡��]����	�0��ׄ���h�E!�`�~��o�O��U0��X��O�ӷ�ëIi۶B�z������Z� �w��G�{J%���I4��p��+0 ��>�ٽ�<�_& �&H
�]�$���w�V	"d�?�B���JP:�ڢ4���qV�ST-� S�%u�7ͤ �� q�#�C�S�Ka3o������|�V��ۋ�X���"�%�(�&��8Eڥ-�ǵ%=��f{r��됚6�[�H
�U�LE�Ƃ�V���Ԃ�Y讴�1%/y��p��Q�[8�x�t�E1�:E���,�H�H��(�F�
�I��r��qI*ue�/�����mC���ljK����e1�*�����C*ų�x�P�Tj~�Y�rS6�8^�C�ے�s��{�n��2��-�GM�WD7袱�@[%��Et���ۙ��=��W& �+��Ih�F�$��S@H~~��/G{i�I��̈����.�,��)���Y!��<�Ԃ�:���ɚ��ă>���祐�)�#Y7nsj(Qw��Z'��"��9hR�Q|���R��_RX��y��,yY���\��;o����4'}<Oz��b��s�X*I@$�0&5!<�Y�����;����ӧe]l�f�0`yI�1�M�ʱy�9��3IJ���yQ0���Np4Q��%z.WA��b��ϴmv�$V��N�yH�Ҭr��È>I�����:�I�lG�}��L~��c�Ե�Uԥ5��by�E��O��J�O�䴓��8Z(0#ө��E�Q�.��σ)�F|��+:��b�x�}����D��(��I�q�稭�YyУ
���jp���U�6��	՞x��Z�Fgea���_u9��ߋ�3�Ǘ;Y�V¯�އ������N��]lٴ	�Q�w�}h�{��
�[߈K�=��%�|�����]��[�Ë�[��÷~��]��h��e/IY9:�;=�#���i��,:Q�J�o�	)
`P����H�e�.aJg&ҳ26E��D�8ڃ7rBRD���>F}��ұ�7p
��w����>�K0�7d���+��,8�*F'�a���H-d����#.`@%;[7mš����S47�M?��xh�C8z򈢱��"L�0�O��	��]��}�� �Τ&����k��,�����0�Mf7����(��C�P�[��r%�h�	�*�3��(�.���Z�(D�(�*cXY^�}���"�NՓn9�H�� ;g���G��4�L5��E�tyu�GG�8����:AO��/��,ϝž�= ����m�L�t�yn����Xf�m7ձ�e0��=gΜ��ɓ@$ۂ���-z)��AM�.��N~_,��tz�t����x�0Ta}�I1X���ҳ���iڍ
Nq�+QbZx��(E�)��v���j̍�<�߾Y���K�J/���AL�-פ�8R����p�kS�Ӗ7} Mh����&Z9��nA �S���A:�*�^�L*�� ���{B��9�ԃh�S�y���<�B��) -םnPض�p�6jP��H��5B�ےO5U����H����-��S�d��m�P�5 �6�)b:�qڡJ�< Uo�\�V�bz���T���>����O��wL��"NX��qpU�L%~����03�����~)�L5v�[����?��z���!��ݻwc�\ý�ދV�G�s13V�/��ǰ{�E�_�+oR��yw������|���v|G�����8��`7��^f��#�pߡ9��ɴ�X[���#��4R�<y��U )VR�(��̥S�!�`=aښ�O.�@��!m����&޷�Tn[�"ämZ�*��ƔӔ����4`m؀��)�بw��"�K�S�HY��|)�^x��q�� [X�;5+��?��_��_��8 �c��X��AWAnJ).�Xe��"Z)odM�\U�(ZuH��L�@E�9���bվ(��4%����M���r�\�/��<�tB+
}-���!n���Xt�ViǴPHSLVk8�o��o���H��)j&m��yO�g/�-�x�����.��l�K4 �sOMjd&b�x#���E[Q��j����ޛ�Þ�YR��O�A�Iߛ���)뺸�m�k�sLr'D�L�ׂ�a��dM�4	�Sǅ�}��tL�-׃�Y+=���)��� l���*i_��SB$��^����ED~3:f� ��z��v��Ҹ�F{~AiG:�����-}f��`X��n����=e/�ɔx%p�b��V`��"-�0P�6e�@� 3�K�[��j~��M��r�	�����!?��PCE��t�k=���l5�@Ӝ�>N��л.�TV�z����=нO�K4 �aT��: �ްv�qR������#.�*�]&�4��u�p���4��SAnz*�S$�DGE@#.h���.���4�2���36͒M��D�U��b������Kn�?����W��0�O���g����������nBӧ�_	[�l�Duw�}/��*���%���~�g�HZ��ꛆ6��7��F<#W`@���m��ߪ�㾇2
�y3�������K�Ҟc8pr)��9�.�!	�G�B�e�3��1K!�m`�� �lA&	��TQ����U:Λ/�B/��/Y=`u�YK2��?b�PLgq�
��� ���wz�dEH0�爔"
{"x㦀٦]�/��K_��.-����"Lf8W�����e�Ey����t��դ��E��ąB�)5����NK�Uzi*���Q6�k��;��7�ԅM�߃/�S���(�P�h%��1���48E]�[V��-6�Y\1W�]���ic��9q4�XT����_���z픐�L�܁��/pť -<v�2U�ʩ�  !%J�0z�;��VX�wb���t��E��H���w"A�V�2�y�n�(�V��:�8��Q�k�Ĕ��@(:"K�;(z��Q��X%-�4(֙���Hݒ%A��>2�����Z4 ����G*h����˟��`��D�+�]��<���H�.E}�I��$��b`<�.��:���.ݽC�<��C!�!�R2k(n�UQ�� ���TBѾ�ѐ�&Ct����R����7V'������Rb���2(�W���8���!����P?. =j����9m�(���z�D��I{�F��1'<��q�Ĉ��q�\뻮q�$����:���(�c(Kp�� A>�o��q��!R�
�$-���xϯ�Ͽ�r����Y�p�e�P��&���-�L|R`rp���u���K�C������R'��6BÂc����+Q+�����F��
fG]���� ���W�h������ٿC ��?��=�����|-+xe��ՙ!`:x�l���1<vzQ�1F��bh?~�m$�"���G�{���w��$�;R����~�1�i�P��)QJ��,�uAG.QJK�� �⸳S��p�5W���9,StNW���R\8�d�t���<��7�F����zSB��ZZ�f�9�]oe��Lb�W�����=S��P�®0�����=PKi{WY����ݔwk��N��������&T)A��=)��8I1U]�?'����˧�;s��a��޽mrY0�����C�S��V�Ugj�6ĕ"���6]w�5����~���]R�T�	� 9`��O����<���<5/i�H�C����R1(`a[E��(���m��9��+�,�S�)�AN���<Ora���r�>�P�դ@�P�S��eP+�e���	d�2J��g��t$�#�5��n_P�f�>�x�-� H"�<sZ�E:��q�Ѭ7��O�)t�f�rY�$�a��VF�Z�]*�+/G��q��`�J�D�)�p��0>�Bu>�B�-'�F�9(�`jw�wO~�����l:(�\�,�E#�_��(����,A��� ��X~~nG��}���2dl!�/�1�	<�
-h�4�b{-�Wۭr;�"��u�Dt�S����H~���q�ak��|71�Q�U��ua��%n��K[h��\�H��|�+��z�P4� �z��g�R��>FN��+���e�W�m�8�L2�{��s��{p=��W����,��{~��Yq<lD1��#����0Q��޻�SM�4����w�ܛq�����W<��a�/���:\��^<��a�+��(��͵�������9 gc-hT�o��v�9�f8� �-�"BLh���Z�<%fWTm#��utu�&!,�TpY��baHv��iK��F��(٩�^7�K6o���"VZ᮳�`����!�i+����<#�T*I����q�U���﹠�mG~ߍ~i?
CNj˅�#�U�]p��qk?Tn7��]��/�K�*
��5g�p�?MQ9%���s�f��ϫ�少Jǜ �������ꋄ���J����\����ڃvi��
+Z�JV��R�L5;�� �.ۍ�g��P�m\{�h/-c߽�����`N��q���Qk Db�S�a�J�m�B0I��B���vcY@	�5v�Y�7W�a������-�X�R#S���<�bI��<{�2���˘�,�������'�
C+er���,U_�7��7mD��@����u�W%(��t��������;��8��Dz��/܊?��? ����C��|�Ա�N��d�%��mL�N��^uNq��Cm0�;�qصqt	@m[Q�4k�����?��jd�s4�QZy^�4@��A  �kI�$kʉ�ЙԖ��49EKylis}����uV׃r��AC�)
)����J6u&l�pŏ��Q���.'%�v[&n���D�׺�;1֐�!F�F ����M<T�n�l����Q-�~�]x��.���@��b6�H�rl~�'�K펜C;��h'�x����K��p|R�+��-4��#���)*��&"�B7�ߵcg�p��=LVm���߆�%8A�}�0�pX@W��]�! �fWn��g�
���z!-��$�9p�>q��5e"�Jt�JȻ�#��w2s����9�*%O�1kAzN����6����l)0r���_�#C�L(4��,-^�ǁ���6lٌz���VS�-�A��h;ʌ�'���ʾؘ��'�� z�*"Xp�"�W*�51��d�H��� Dk=X��N�.\�N��>ky.zL_+�4���vd-�l-�-*\#vy����)_���.Hi&bn�J;�ʾ�ĂJK
)6�So!�d�A��4PT#iN�L�.B2�-��6\u��!)AI�k.}�F��{?,=e�9��3��@9X\s}��<vr�)E}�d[���=SgF,2W4���U	�t\�1Qo�e�啊�,�ŝ*�dr�CJ��5j�ڢ�ँ��p�n����gt0D�M�W����,��^�-*��zXYY��,]����Nq���8�x�N�P���|�-���~�����<��󝿂������-|�CS'�?�F�A � ���Q���(�N#�<4[<[8��Nܩ	��txlW(c*�n�@�?���R�Y���9mK�L�$���=u}H !����q�
w{�����I��N�P�^	����H����ߓ�ɾ1��pKH8Za.M��-�_]A���S<�����$D]���$
�Q3TP��^��n�Q�0��i�UP�L��q_���Y�2,ҿ������o�l�1�E_�'�$�:m��9�a�-,ԥyR����h{W���l�VE�-H,�ǩ��hu{ط� >qs-��[D�XE©'8��c�vL�Fq�]�(-M`z��_�ŷc�ۯ��7\5������p��9���    IDAT+0�x��<��g�
<x�P����(C �	�]��⮃�����L@H�^f=�-��j�2��;��"LV�P��{�Q����i��3�S�T*���ԙ
�����u����[S)�"��0���谄�>(KWq|"�+Sŭ��	��(V���I��N�_v,�)����;�P�X��-<&M��L�-E��{:���6��}n�٧����?9@�ɵ�K4�
&@�c�����3]���$�W.E��8eGU�1Sq���<"�A]E�:S�ną� �|}e"�(z�v�k-Bt�Q�`��K��.��Q���{:��x��w�PԓO�.�]�����x*{F�ʫ�Px���>�6�9D�VB�D�N��"��j�
~�ZU�-�__�T�h4�j��i6��LM�g����f�����
�-�d����*�� ��6)�a��j�rYrT�!�k����~jjqJ�
���V�c��V�[D~�?����/�9}6{�{ރc'N�kbrZ���~	� p*W+�H����VA��IL���F[�@R	<���k�6��Xْ��hit�[j�.>ϟ�6��H�H��e
q�o���Uơ�������rG��L^�u��,Q�r�8POל��tVY�Z������$��������'��ٷ��]�o�>�U�����B��Ut�#��)��İaWFs�(�/�I�Lw�{#��"��!��������	��^ZZ���T�#��j8}�4N�8&�#s�Z����Ԫ�#��@&�6N��+�v�G�цaz0�刞�*�"�qvn߆�� � #�03Z�{���<VB����_pŰ�z��݇���Ë�;����u~�ɬ�G�ٱ�cO��=����9�c�=ĩ�85� Du��H�Q�XU�j��$"jME +$;n�qS��|� 7�K���$�B��kv�B��ߧ��D{�N���0�H���
��q���sP�2����%D:��ʨ����%h�:�^�)�v(�s�r  ��Z�0�s;& t���7�U3�D��eK!��nA��I}��}�W	��E��t����5�2h�*�F:A�S�p,�ǯ_�j}���6��(,�sR�( ϋJ퍛S^ٸ6F6�G�d׷'��^�\�V�x�{�8��r5ʝ���ֱ*��*�<�tL��I���i;�*ӂ���x�6�����ص}N�:���yW�%���>�я�.�%�s���{���e�S���$VWW���s����{��j��������7���l|����=�䓨���+�1??�O|���\���Y�8qw��_���ؾ}+���0�0�;��y��*F�%�m�
���[��o|���������8z�8:>�Uj\R�Q��{������{���?���Q,�����S�� �?����̢N;�uQ�3�	�8hA�2c�TH��Y��tr����>�=A X *�3?���|����űC�!
u=����OJ3�s���TQ@��&�vT��-?�T�2*����cԪU��0������<�*�R`�n�h��S�N�-	e�S�0�[���.5".ܱYD����98��#��<�*�o�pi�L�c��	tx#د�M �"�_�o�k����uZjZa�d!d����p��T����� u)4;�G���L#���\��W�}�ܫ(���9x�O�	[FK��e���]��]o��F���<��p���W��}�g13�+�|pd����^�\������Ѕ��5# D
A��.8�0����5�1b��j)*X�7Q����:�{�n�n7�$�p�а`
�dp�.+�ۂ9R�U.!��*B%�����ȶ�gq��ZI/@���h!� Y�OT�4�\�m�WPTt'E3�v��z^>����aw|n?o@�`r-)s\�̜ҥ��P�.���Lt�^�Կ~���d�#ek���S̬����%A0s�A�����H�(�Y��(Ed���Ǻ����<6�V�S��a�-�6`��:�<r'[ꋸb^�:O~�Ŝ��y<DL�h9z^&u
�i9ˏ����m�o�q�Ћ/5:|*{����-�T��?����9���K�z�׀�������{�W�?������2��~<p��8~�8V��6� L���7~oz��ƑsK;�<� Z�6�:}
?��� L�Lc~~�`rtL&sssB�9u�4{��}����u�\�������M���7^89z<��]_�G��2����8u�4�O=e]\�vL���:�1\����X:?�cG���O�K��&���.����lAZ�olvei����A�O{W-��G>����&!�����a��J�|��X���v�B�qp��_P��Z�.�� ���yj�����U�C^+*�T�L����J����i�{�5W�K��G��T�:�/7� �fӀ^r}���B�����(Ck�x���6!2=D��^��bU�#i>�d�=�������ò=�����S��Nj3e�m�(� !Q������dR��TL������!�O���o{�^��܅��	<p�T��>Us��?�&올(
֍Wk������kV`x�|���~#+p���d~��umt�X(O��_z�	�ЂY�d2@{I���!n"�V���{S�9�h��U�;���L����Ba�:;�,�h˚��R([K�)���.yj�@TҰة/p�LqU���I���J|&�$s����#ȭ���`1��2I�.��V�"�v��zF`BВgv[uVD��r H@���@'v������+�+)+-��b�>��nUyr����\@��+��3���NUX�ֹb�KA�ł�BF
�ŉ�<\�Qz�&ǀ�Y)���r	$h��h(^��X�NS�7�](�H���1TKe�	�>uJ�I	 U"mZ��L�<gE�L��)0H�R
V,z����+�㝿p^y�����l�އ��ZG����}{q��)��60>>.�R�~�w~W��6n����Ç�����=8��cXi712:*�^������<ﹴs�����p��:�$�<�O&,=������136�m�����,������}J�'u�l9��~�=�y_w����)��?�,,,Hb9�a:p}��e�;����)g����e�l6��)��H)"��(� pū"^�k��yA�(�%$����l�M��l;��̙�y�s6����z-|{x��2�3���{�S�Ⱥ��4j}�)���x�ɧ�{�N��8��$H�dd
��� [��j����[ĜB3�dr���I�*�I��b�J1\O�_���Oh����+*}�_ �nCE���=3���O��*�=���W��)��a�lrԆ�jҡ��d:�N$d�JClD:���_����ú����Ups)��ǩ�⹬�5��G����t�Z�����n���Ha���KѴ똂���kC����|*�&���-u趭h|�> ��---hnhD]}B�_�l�t��[И��q�ݹ�6nF]K2E���D�R�fED}�j��}2,�O�I����`ތh�k��e+e�h2�5�+?�~L����8�ȉ�O��N<gb��
L\<���
�b�x~�$��#N�@�����c�`n%��D��@T�YQs��t���� ]&`A���G�rE����S \}/N>c�%�E���h�\��4g�E��t��A��;99�,��WhVW�Jb ��u	ч��l<��`Uq9-P-j�y89R����#r�pR��:S:��Q�PF��
@�"E ��C}����Qs۩N.9I�T5 U{�U���rB��i�9U��+�R�vWr*8ղTN��i*�������Xx�}g`a�Z�h��4u��g`h@�=	�s�Y���)��nӻq�P�*Œ��H�W-,��©��ݨ��*����Կ�y(@����LMAuX���C��рmu��l��x�Ǳn�z��K��Z��~��2�y�i�j��v������}X��
��ۅD}��Z�@ _��z�L����r�7l��ܬX�Ͽ�D��H4
��Y���~���z����/^��߾s���?<�6n�$�$U:,2�}÷p��_u�����z�ع�O^���󟿔����.y��yο��;�9I�	=X�|��P�����&�W�:����&�ʮ89��G�h������d�j�\;=�uM�絚����D{$�"�� �
�ٜ��Ս�i�����%�~)��H�u-�=�c�N@���hc���UM$i�m��@!W��llE8�O3�Mgp�����ҋ(�#

03��6��l?�<!; S��B�����I���E��d8Z���Rʔ/���CMW�\�W�UqPʌ��7��s�z�h��uEdp�!���(�[��BX�� ����X�r��7C�
�_��3:
���D��G����� <̝1M�,{a�P[M���Q���#h�}��A�s�k���X��t& �_�r�{M��SKV��\^Č,�S%kwቕ�ظg�E�Q6�"p��_U[�����0�!`�4�T'N7Z�K����`j%����/K�A4h#
"�#�N��"C�S� \�2�0,VC���%�E�|� �wTRrX��H� i���v,
� �	�d���U�+�8W��#I���w{Ѩk"�V�wU =nXU�I(Dp����J@@��(U�)���>�F�Or��uk�I9�~��b��PM���p�t���$������ۍ�LRV,Hމ��$��@2�bp3�����$#� �lnFCk3̾��J�
�HR�9͢�o �D<����ZA<}���g~)m,<�h%T|2�H!!�E��۩��I�Y��uw�9tL��	G���g��p�Ņo9u��m�~�w>�E�c�޽B��,[�Ûn�Q�u�?� ��G���}�Y�ٿ���3D��6\��/�.Ñ����,�W�Y�{~�d29#a�!���}�K�li��:�*��]x��'���Ų6ԥ�45�+_�7}��Wݿ�}�y��o|]�3,f���&^\���n޾ݿ���ܢE�N���(V,� �ijs�.n�j�<�� ���^��\W�V>���\�\?W�?D/���+����� R�0w�4�&��8e�q��	߅��LPK���s�t+�������4^�T�
J���`ŚZ��D(P5of�,_�\rT5'�l(�Q��xB�R��:TܲҼ��)�L��gx*'IV��I(i� O�Ph���+ߗe�[�`!��8�%F�aZG#.���q��'!P�*s̈�O=v�K~w�ֶ;��q� .��'+�DK'���0r�F4u1A��38��Ϋ&��;s�uX�t��X���z����h�2Cx�^7QC�&+����[�����X����Y�^��ӎS
b�B��aM�<�R6��� j!XDHP\��_�˫��4�q�w�r^�Y�>�\E]4�����]F"l����S��)N|(k�
o�r�,:2YeGǾ�I�
V:ȗ�B�g��4�,\�i�4�
$V/,W1TU��e!�bS@���)T�����[+�bʹj|�Q�1Iq�	EU�.�rZ���4`��:�U�T�[hM�\�%j��{0���^�������I�ψn䠐��|�q K�x�*�.���x4�2)+���CpW
6��JpR��>�<�5��� � ��́nD#�$�J�.Z�x����t!�a0�Lu��tMÊ�/ ;2�~dHG���(���*D�M�x�T�^���P��s���;^~�y�[�����{{z{{eI,#���:��{���zy����6l���>�ͽ[am��i̞9W^z9u8�9��f������5$Sɟ���L[���S8�u�a������}G���X�|�,��!����Yo:Y�������O:N�����e��t���C��^�|��u/������`�}"��:J�O� W4�4��H�@�jhFNҺ�w�^8~.��k��*w����K�����'h�D�_�&�V�d�jB�6�841؝��:�Tl��y�}@0����_�R���P��=��szf�C*�ACc=r�!�w��e��0�n\��*,R6Mt%�p���j%!��<��Q4T�;�$�
 ��! �yK2�}1�;���{�2Xɥ0�4����bR#� �L��cfcB����_�G �M�ڶ�_(���a�n���{�p�X�z�V0�\�$ۢx��L��x������cެو�X�d�L~l��>��cZ������O�����'6�n& �?�!�ؠ��
�ܰE ����& ��۰y_R(X�s{��r��eD�;5����h)��/�a�7���0��hm�B+�Qo��,�Kd#�L#"h���f��?�[�`��8q�C2��0��"+@�E��
�7We�K�$vCٵѲ�|���!S�&���'Է���`A�R�U�yu� �ve�)5�;T�!�q�t�����)k�?ƑgE�C�H���������j1�
�q�2��0�E��s�3}�P�!�x�9�)^���<m�˹l�HX��c����&��J0̉!���	��XӦ!�KcP���+���cQ�<fw��*R��8���0� {w�@�t,�,i�^��6Hh�R�rux�إ���9 S��{���8z�4�s�	��5|�]o;��xՋ�t֮]/+)a|�����#_�y�̳���?� {�I$��RO�#} �Ϙ����kV���_��+�Q�d����ÿ]w=�9���ߞ�Y�3��w=�/��.?m�ٽ�ԧ>����<�������p��Gh�=����}E&,�HH�8���x��_u�ۺc�����۶oǺu됥�ʌ�Ac�2�
������F'��& F��}�)��z���Q9b��Id�
(�5�\�n):"#kV�r��C2]GΕy�{�,~�)��t�m �Ԗq2Q���H�F*=$���E]'���Q?�
��@�T)6'0�ϟ���<�=c�$�(�ߋ�}�K(rB� ��}f�%���pF�r�R��a����Z��6���X�g�'��Z81�ꦼ7'�F��!���w4h@/�q�މ�.:( ~��\��V��c��)ǧ�i�1���X?���g�cኵ�6���P���C.�^"��aT!��ļY�ű�r=GB�#&�p�G�U�^Ù�W����X�?&.�?�&^�^��k6
K�b��i&^�9(�-�i�=K��Y8J��x�W;�U+u'#�,��H�ES�����eaV
�e4EL̙5񈍺�(b��eM��H��r���e��ً�-A&�2*K�Ŏ��0>[���H��HH�{��(�U�K�����#š�ɦ5&���T�J�����C �I�08����I���s��K�_�������J�^�;�@GUi�NY@�<z�)V_U�\���_��hH �u�_�}��\����t/�|V�"B�ᴦ
T$;���Cww���H��B�����{Z�fd�H�R���L��D=m�(y�e7;Ă�XD��L�/���hg�<�]aI7MD�A������;�0�w�|^%�3%���`�>�i�Fq��dWYN���}̝ފ��u6c\p����޼���w���[^@F+f���q�mX0��i�ǲ�����xf�"ttNB�X��{.xN:���C��<��5W!����"a$G��~���;��	��e~���o�{����	ÃdRw�G>���>3�N�x�!��*��Ww�_��W�X_/BwR�[[���s��ٰe{���Ïb��X�b���`*zc)���Hб)P�p"ǹz���8r�!	���(�ȝ��v�U핡 �L	�E��	�k|�������鈚&�PL�i*/��Q>�\D(@(�c��ǯd�*6����ـ x��*N8�D�w�۰c�n��)S'��+�p��    IDAT����һ~�A�4b ���2����W(�P�ʟ�^Gɡ��S�<�V,����h
p�k�@�j5.��Ju!M���}�Lm4�d2p�%̝ܬ���G.��޷KL����X�E�{���A��
��/ێo������P1�Us�:�B��'���3��p>/�s(���.�뮺�1���	�k��ص���  ��k<�	�D+�$t��Ž�ɸ�)���^-"t�bS��
��|��$U�L	X��J.���fGP�v5bvgza�'�p��.Lj�C,d��>�bn�ܘ�<+!oP�!�[�D�jLv�+zw����f��H!��mF��ؓĞ$
�߰��,�)�F�D�UꁸPU����Ie��sJ+Xr���}c��.��,p¡�j�UA%�v�E�}(�D��U{PWr��R��B�&�ew��	Iu����V��GI��y�j����8Gi��j�S��T�(�Q�:�Z�����P���*N^ҩ]v��i���5&���e�u�T���+�i�B<��i��$����s=Xuq���%厇��	�8���b�u�F�ߵGt 5�#v�%�Dhc����I�<���2ݏ��"�
��x�9o�_N<�0mӦ��jq�v�f���(�$��mC+�{��;&r�زe�O�����C�߲YB�jE�uĜy���O��k�!�y��'�/\�E)T�A��!Ķ�k^u/ڴa�����=xq�j !�Na��n|�ӟƩ'��=�ܳ~gg'f��Ю��Z��'��DG�(��'��ox�!��q��g?�Ml��E�	b%���F�ex.�K>LZ)k��,��y=��& ��NjzXb>�@�<����<gV�Iץ�8 ���$n�aj@�K�_gwMC�0��g��J���({�"Ah��7��DL�j���Pȥ�J�aߞ]�옄��QD"9��=s�	���g��P(�];v��t�ǜ�f!�M��*[���	;ƾ}�d����*��o@4��=�0<6������hh��b�D2�����F�XD;:Q��!N�!Nyk��hZ9�������Z�q�TI=_�m���摢��|#�<��X� r���02�$q>z�����h�F�>��P����n�?��6 oDd:�9���Zʉ�@��`���騋$��������>{ه�������Cϩ�[�ĦN���}& ���Ll�?�
pB7	�򁜯a�����5�>�����m+Z�$]�q�j���5ȟJ]-6Z�@{�������pfv6 a�H���M|ǎm�dF�Ɍ����B�+�iH��-At�zf��s
��z��:�����;��U`'�P��10Z�H�{�sB�)T�5)R7�Zs��G=y�5;^�2����~Jb;�$S���	x�W��M1�~񃪀�:	Q���C&� @vE�6ƅ��BD�v4q�H� K�j�3ߓ��}F�pD��
q�hq�� �
� �y^�)T-_ϐ�_��}%�U��bO�	:io\&�u���$��N�3
|:*1p��
�ts9�x��e�vP9iQ������#p�ydYh�O`Rk;�q���'�6G�{Tǝ�K�X4p��9aH"�2��Չ\"��3&�7���z����i�w�_�҄�S��y[/n��7D��J����|�t��r�X�v��r�J<��cظmB��l+��Sތo|�����/��8Fٕ����׿�M��
����y>��ً��7��^�Ҫ�>�ۿ}�شib� H���(���
���wh���9o=[[�n��u_��ry��僂�k�����JN߾g�OpB��*��LE��F=�t�"K\q*0lfV ��X�ȳh�l��{׭����S��皶L�$Q~��W��Zn�L�h=>�S��e�K��	�YS�65,}�9x�N��t��],�0<�v^x�Y�3{
���B���-!
c֬�hmj���D"1�����$�c(��8���#�����	G�q?��DX�Ѩ�!%q�§��wK�J�~*��e��Q�Q����"<�e���i� �Ew9Z�C6t'��^č_�,^7w*�B^������>�n�̓p�L��uj��:��Z���O>����V��x"�{�����=H#����Ġ8 �P ���B+��=�M�x��g(r2�9�+>�^L
y��q��'M�P�H7��m��Z�����pMl���
,^��/��bhȗK+9�>��C�6a˾r��Xp*�h�D�7đA)�B�2ր�p��N8|N9�0tw�a���л~���@{�7�(J�<��
3B�
lSQk$3����I��J">��5g�����=$��w�c�K/��}:�F���06o߇��
ZX�t�5]�l�{K�+ "XBuv�ԧ�.�9t��z̕%=X�ۮ�pS�hjlA��©�TM@�'@�79�=8=Q�Vv?%՝��Śi��$�2,�A��.�Qt��i�vXTW�-w����P֣
$Q*/,3�Eze�.OҾ��L1��@��o����8��v�nY�P�!N)ʥq�U�.��1����z����2Jt r�)x-;�褓�l�P����D�0�H�e���IF{S�������d 	#36*+ng�2�����J�B]N@�0wz'fMi������w�����+Db	����q'b����}�F��y睇���=�_<�h�_.�<������޷V��mm��#hki�g�����ݿ�����)���cO�W_���3e��h��?��p¡���?����K��S�c49�PȖ)���
��k��'.�\�뮻����_�:(�gw��~�L������%�n��f����{���yk�6�%%��S*� `�r�D���F��`��p5�X���@�p�lF�z�C(����(��5�X���T5�C�%�	�F0TV��AP�?2�rq��y D}��Ć�*��$p	�h�É���Yo>�S;�\_'�&ݗ�HDc�; ���&�*-�	��̙�Gj6�|����?�.]�5k�!_�o���l�ix��%5�Q�a[�Q"5����bs��^�`�7u �����~��=���z�6����M(�SR��dm�124��x�\��fNi��;o�6�d���1�G����}�oQ
�1���R��S�W�5�<T<~��7g.Z�[�h���0�5��.� 3��p�p�)��`�1�+���������+^�+�h�q Rp�Ⱥ>v������n�p���݈z�w�|zݓ۰g�f�"�Ϛ��D�V���|&Mj�ε/�G����j�i)fe�\�)`yc����&�Cf@C�)���A:�C�))0[[�1��h�9CR�����6 c ���L�6�I�W���0B��3�ʢW�ﯴ�O6V�u6�I�ډ�!�C�L�i4N����6D�Kg$�0�M	����!��L̓�)
��GP,����t��!�y)[מ�VF�+��Ej҃j"c�(��0Fg2�<�%���sh�iJ���	���HHR�m�F���B?s��9&�gL�GM��@:<v�	>��؇��y5|����M@�L���(��)�V�+}?B�rɢI��� 
��Ĵ,)�)4�È�C�RFW����)�0���X�dãIDc	�$����9ݓ1��{�o�	G��;�;�=����m�����!��Kw� ������8�p�UW1O����� �<���^���(�024,S��.�8>s�گ~�k����L�x7�r3zw�DCS�LAh9}���ԎN>g�����b��]ذy�lX�\>
�)�&أ��\�K/��v��7�3g���f�,Z�H�y~q-�N�*S��3�r��(�sE<����P4�0�ɗ���J�.p�D�D:S@�!�
(�1���cxd�p�L*+�#b����Ȥ�0�P|,���:򥼲N�j���|(T^���+A� <�u�g�DXױ�A� ��E��[���&�����M�fF�,��R1����iSE|޿{��k����݃YsgIz����E5�o��~�R�Z�
��2�4Oǁ��$L)��#���0��f8t��t��Rm)h�҄T*Ex�̛ކ�~�˨�=�=�M!��v�7��V�-�(����]^�aѤ4$�WJpJ��K�X�؝(g�Ќ0_��|�g��d���% ��·$���A3��ܙ���8	�.�	P�҄�x�/ČfHᬓ�-��o��6�����l��[1�+��Ͽ��/8)f	@
���Cy<��F��>���OJ��{�"�99����H�ߎD��Q�bAO#�p�ǵ�ޅ���+�u�Lj��Y� �N!�P�
6ǋJ?�n��#d���JJ��4*.� ;������b��݈7����G��-���w�?	ݪG���R/n�C�"�+�Xpa�����읂4\U��Ң�`��af̝P9ܶ@8�ݹ
)(fy��R���o�(;%UH��b6�i������E8kl��{O���2a�F��Ja2mU�:tKW�jD]���\X� JEI���U;N9�W�1�fx�� �L��$^R�l�W��Q3�K�|S �o�$gP�_�(��r�ID�0�
����e2B)��n-#�\~�łS����ņ5�
��B�r
Y)���ϑ��H���9��ք��)b�ڷc'��K�DZ�C���mh��at`7�v֛q��Yؼq�L@��ۏ�/���X�5/a ��4������y������GC�&�ؼe� XN�!�TB�X�Y�����>7l�,���{a�xv�"��S�9{�LN@i��ڎG����.ҹ�d��ܻM;	@,MC1���|������ތ�K����]@���_�2+N�a�	��>f�P���ի���&e��_�h�\�rN�C0��HR����tC�ď�!hG嘜r�)8��s���ŝ�܋���pBN!3�[��ޮJ5d@��
A~-@T4<�B[�湨��5̙҅�e) �l]M$�.g'�^'7z�����.b�b� �O$�u,��b`� ��r�,F�#hll�{.<�T���_���ݼy#����?Y���)2$��`m��ã��?�:��!����|'���8n��h�� ����+7݊��ȸL�7`����v��ԇ5D�,����v�����7�����7�X3ʚ+���Ϛ����	 ��ҁ93f����/C���
��܈O\�vt7��Gp��sq�Ana�1��4+�?�����ˉ�X�?q�:��碤��ҟ��K )B%W� 26�<��&*���0wZfMI���;q�aX��Y��������7u�,Z��A�b[�:�������?sAd�P*!����ԈPJ\�l��$3gK>z����?�y�Q<����uƦ����������2%�٫�n�֠�����G�i(�$,��y�!$|��]�f�=\��c�,J��$[�(��s:]�|�&)�%�4>ljhJ�G��]wN&4Mm�����M��iqr���1�(���i
��4)V%;�*lUi���� p���A?^d��5U���#�P�D��O�O�mbP�hw���`HM�jnc|�;���K��t��WM��lՄE�X�����?\�I��`���F�-Lio�	�sg��.������. +�ͣ@��
��Ϡ!���4<̜6��q��iik#ɔ�A&���a)�u6��1����׬E,���hj��,�Y�P��475�1^�$5M�M%�'%J�a��)�	$�q�G�6y� 	��\��#�I%e���h��W��"axm��඲ �ߜ�p����d��3n+��g�өg��EHqB�jj���ס�H(�t���� p�+'J�fc��FH�4����߼�cڋÎ����ǞZ;R���!�(za�R�Ft�BX�[(W�-ޑk4,���d�L��D��R���5 <ߨ���d��7��N?	o>�X��n��߷��W����N>�$��9h�\��ܹc؟�ݤ-_�ַ��G���[n���6lX��Lf��d<$�Ex�[�a���o[(W<�na�'�����	ꨔ���+��׮CO[#�b�&�i��������\A�I�@ǲl+*�Ssaz����cm���?��A[�=��/!���RV&|�8���$�,�؜��hij��V�X����n��?p���Q�y��j�mf�i+0����N,��
L� ���6�٢>;���l���#�^�K;����7P)���RQxh0r��q�QS�=X��o�ُ��dm���B��kÊ"W�%�bT�*m�"��X4"n6�YȲ��$ba)r����X1�ypl��'`$���n���w!�Eџr0�r1�qUȚg��&�s��z�@VܥȤ��pJa��+`hl�@&9�p<"N8S���=p&W�p�@$$��t� W������-,qv
h(�h����pri>bѰ;(�6�A��I�1��[�	��XZ
e�n@lÂ�2���N7TaA�A���^)ò8�V�AS�E�"����RQ��	�L���;��d���:թ|( "�hʊ+�,%c&�
�\�jYt]
S�r���b���%�A�#��Rv�@.�c�bRK,]����ػs�����׶�sٲi�j��DL��(���P̧�����e�py�XԖ�H$���I�Q_� ?/��#Ud�M�1<<����
�����ۻM�hioC6�C�6�|o�C<13����h�H��6��`g28�߱t
�P��k��М F�������6�iY<8�@sk� Q>�6�u��t&#Ȝ�j`Ǟ,��/b[��H��{�%�0c�|����s�iW~�V����V�Q4%>E�<$��i�Wr
Bm�zߚ}�L"YUs�� M�ԩI��X��@مE�j��H���Bn�{8�~�i���������;�zq�1G��k� K�!��@�_Z!�̻��Iɏ~t����ѷg'�����a8]��XFM@� ~߄uN�G�sjft%�WQ \��H 7<��+p��n�<��zzn��gp�+!���4�r�ƣQԅ�Y$�.��¼�:ma_�?��+�E��� M~�p>*�}�f���w`�fL�F[S;�-}e�G(hb�N\���t(��-�Νh�NT+������.���^�+�l�&@4�1hZ�R�><�j'���k��*�dլ4Q�%*�p���ⴣ&��7�CT��eO`�o����KW-V(,E3�ϩL��vL뙇��Db���7�ݚ��V)���TC��X�d��QDl�P u!^AhH4X*���,Z:����^��1߿�N��r-d�0�2.�KH�	2l�D��&�|��ՅrPb��
�N���4<u�7�{�/��l��H(��_��EZ|z��>��~�+ؾFs'��(����8����S��Ɲ���1�'P��R�E� �[̇����\ȕ�m��a,��S�.�CxN�TL衸P�J,jMҿ8?�q�<B0ڏƩ�����NVzذ~7~��_`ժ�Z��J&Y/f,����h[�^+�b��q�0D%*�M�����ے2O����%�Wv�j�9	sk��i�~j|�5�ż ����!o<�8��t���A�	���d��1X1U0Qq���ɇG�[�݌�ځ�P%���L����m8���D������Ϝ�P�P��Dc1�ҕW&�7�S&z9���Yd+�Ek���pi��Txa�Yr����u`� %�L��d٢3�[?/Ry�6���DDM)՚�w����&��FRt�S�Ϫ����e�ha2	�B��+�X�����o�P�"X�nn��W���Î�@�!)p�æ�
��R��ɩX�E��@���9�VH�0g�t��`=��
��S�,*^��t.z����3O����{�������k6l�.z
�b���3�M�v�{w���Μ�5    IDATN���J���e��^���	4I�]%v "1�'u�LS
0Q�߅<�M5!�<M��G[�Ən��1hSm��K��_ݍ�na��-ǅa�����x$.d/��"�g��]?�^r1+����{���X�T�B�ښ`�|	�L�x���}��v����S��ډ�KVH�{�`��I���X�1�y� ymV{��X�?�K�o�1�1��X��e?�/5�@���xq�<�n/����ۼmR4 E^�TFC���p����W.�@��%�߱i9��|jIf(���#Z�$��X��M��}���u8�e��n�r؇�h�$Y�$8Ō8���R�"�9�,8�<<��J��P��P��1�ӱ��;Ga�Q���*�"m�jV�pӉ��H�C.�Θ��/��<�(�w 뛺�����e`�g��.��<,��Qm��O�?����/����.�N��"X�6RL��{n���j���}�kv�ږ�4��(�¿����%���e��w~��4�[�`�o�Jx��U��Z0A5�4����'��FV�`��* ������ô�J�B�>��j���Mn|x$<�jJ<�d�K�!g""R�]�@-��~�\��2M�
�x���ŨS��8�.�S�_��T�.nK8��?K�{
c�"l����f`�X����f��f�B���m�)�b���S�s�o��j�6�X\O�v�qP��@$��o,%�gAN!smjB�!E�6�U=OhPL��~q�`�m�|Y�H@��c��굮�n���G�Txp�D�T38�$C�Ӫ.n\?��g-��A�:������։TJ�I�����l_Y.��,���T���B����M\@λ�B��3�_�}?�{�q A$�$�:�|�$��)9�j�ʉI�`̀�]+�is*���̃Vv�b�B ���z�@�e���p�����w��-x���I�)���]�{�_�v%\�����	ܽ�c#I$b�\��HL�r��(����_�;�{�tR�\�my@4�X{
d7|��
˔) �)�(e��Z�~��h��c����س���{�3C��3���/�nK>J�-���k<r����� �{�Y���a&��w��0��s�9%�jVT������nt6��痣R�e�;sj+.��h���$�xݼ��:�)�b�9+�ZZ����t4'����6o��2Y���p��`+���s�`ն~\�M5�gGU�~3�<|�_>����6/��_���
��BuȔ}X�&�L����vL�:�ğ�!�l�7ox	[��CzhgT�L�R����Ǒ��/Wp�;.F�����^�j�k�H��XV�K�� `'ƻ�R�H�D5��ŘG�`��f\���q����+�i}cy�R,
_���I�Cv�/�:�{��i��?��E~�ܦ����'x��hlC:Wߊ���݁������{��������#T�`VG��}x��%�l���~�{����f at��U���i
�K�c~A�D!=���u~��+����3Z�ن9'}�߱� �;�+�D�� 6�T�q�"b ]y�MQ�+"�Y+2�8H�2}C�K*3�	Ѵ֭u�	L��R��:�����*w���+�������Z���(�����](e�$0�-ED�����M�����Zid
)�:7�X�f�E���LV��fsjB@��PvH�
�=tM�63�`�X>�a0[�־�8p�AJ��8)��TU�P�I�A�NN�:�e�B��\W��}����.�Uk�8��R�2A��r}r���B�P����k����(l�L��|O^s<$�\W^u�8�\T� x�)��~*�ʊf��n9�lk\X� C$����͉W9v1�.l��-��9��#��`�ҥ@.ύ�Z�ӫ��APY��YSqƩ���O~��^S�[��=3g��M}�(cڌWk@�N���7���lĮ��0s�l��MAȮ�T�e`ۜN�B��.��H
-]�cպ�ȕ\�C	��!�`�x��Vx*S�Q�r��	Y(��0�1�}�Kh��I����q�/~�$�~0,�T&���	
& ^�W�s���Ll�=�w_r5<3���^Qp}K��Le��8]tJ2�<l�4Ś���K�Xq�{&7��#�#�pڱ �|ӝx��oW`��{�'v�����u|r�	@H��C�xy
X����#_1�U�E+�Dh4�X�e⾛����-��}�.x�Q��S����� 3?�=s0y���W���ݽ;�����A@w��ڂPЂ���f������8���O]��)7�6c$gb��]�P���4�Igw�\zG�O��}��߃;�~���n�?�S=���$⿮庾=���5Y^�n_�?����5��0�;�b!����ܺ�ԫ���؟"[=q�o0�w����z�ݱ�?��C������[��C��NIG�*����S�I:��y6����n`�r�uW�o#t��~z�3�~t���F��E(/#�cb]���<ݷԔ�e��5��N
t�T����]v�<x
�`�l��Y�r�!�M�2�Q�K�/-bQ�C'���r�D�M	��$����&��KR�'<wẛ*��Y/R<�>X�X���8.20R4&�{X�ST.S	Z�
�6�mXAK���~�<��}8U���;�]9� � �X|r2�������5��^U�4&e���Ő9O��TAץ�x���M��=B�b���2f�Z���pJ���ru�q3�)V�Ca:�&�zU �A6��%�^����9��Fs�إW�o� r�x���qJ�ʖ��'�˴C��B���jr��7��؝��S��Nc�֭���dJ�r�'�L@75!��G.��]�W]/�������Z�m�� 9@ƿ�C�Ib��h�4�U����_�_|i9���)3y�46t �%������'���_F߾A�f=�G�i���B.SD��
!2i����� �Jp��W8�0�Sh����W>�9�-�\�[�ڢ�{���z�{w��өЅ�'mtI�bL��/��(�
����O\�U}���@�T��4�z4�u`$�B�Y3f�.\�e/��co�;�2��,��������]wb&V��
��E��"N��kq��[���L�uQr}�V�����X�s�2��
��Sʡ���+㘩:~��ok����0���b�pE����umx���}���Q�����ӏߏ�h?�cchok@��AggF�)d��������kP6�`�w!]�`��1�eXH�ub)�yՊVL��.`Y����o����g ��	����#))(�Cضe+�vGq4�!�##X0]M56���u���7�?��(����2X���ߠi���3:NB��]���Զ}N���i�g��۶g��6�w4j��г���|	N��v�L�D\Dޥr�RA��>t�y���C������݈z�LF "֩ӗA��>�r���YU��>�c��	�ޝ��:E����TC�����S��+*V�x��>�N�"�tZ�m`R[#"a��Bvl(g�Y�:����[�&ĮU�.5]���߅�!ES򔭱�M�VED�U�cn;5�_	�	�s��(@�2���,��M�V�>Q��ߑ�şK��i�d����xB~OA:�E�O Y��e�4��l���zYժ�k��T]媀��WF��V'S>G�\�s ��zN�؅�t��D�sX����Z����YÅ�~���(�Y#��]�q��D!�@�� GI-#�1��pBE�8���ìK@�$��J3�B*�d�d�h�2����00���r^~�^�q|����޾��g���<u��}���!&����z)47�
i��S�i��c���b�K�L�45O���y�v�ް�t���vnڴ�Cc(�1��J.r�l#,�07��Ԃ2�X(� =8�c"<� �p ��A4�����0�g2�cC8f�$����|������T�  � uA������[m�������򾿫?�T.�l&-E#�wo���GP�#$(qb��;�p�F+��(����%���ߎ�%�ӎ=|��z-��7Y����o���ϲ��o���� �� ���Vn��=c2� 0a�Y��:�j��������%ܾuQ���{�&�-�hhnCϼ�:✿�5�;��ܷ�6����˅�u��3E#B����V��O]�5|��k�w��@��IY�}{�(WKe���� D��н<ʅ1����n.�v��m��O<�ã#[�8$��3LJ��>���=x�)�v;�=��#kEɣ����|�Z����TS���9ժx�O�w�N��5�恅�];��<�M'����]����7�_��0����Vh�Jצ6�W_y9>t֟/������V��������;�>��PQzw�"f�s*�Z����)�ŢRx�榀Ǹ�D���~�����:"ҝ� S���(:��IA�ȼw��2��2l����� ����|�(�'�ldHYժ�x�p\>/��n!_�ɇ����#��5�<4�!�մ�5��fQ��Q�|�jX2�F���m)�I�b�T*N8�R��W�N4*����I�-V�
\$�&x5=
߃�1>G���)�jq�3�>y��hU]��惹�հ�w���I!]3�p$������x=zw���~�c<��B��z$�He�F��2����q}qW��s9�ɫ�E���=lX����pF�2����+Q�c
��4�Q��B���.A]�D_�v	G��q�8�����a%~��&��ј0�FaV�dJ����
��BumX�j36mݏXb2Z&MC��`,���H��ͨ��c��|d�yW�2�+9(°Z:�T��b�M !�bP��Q)�o�Ɨ��Qo�(��4r��ɇ��H��05S�pj�@C�'5�I���',��S,6Xt<����p������1�뛅���3=�U+V���^���.��;��4N?�����g��Ml��
�=V�V�=6~�3'V௽+6l���<�$��J`Ŗ�xj�l�=��'�-n%;�96���y���cp��n@S�G�P��2�� |3���YG�-��W���V���lZ��z7�Ҋhi��"u��O�Ǯ�,~�1���{k���by�;���)�({��3�CY�Z��C����-ϋ�T���ug?����dF��F���bcI���C�]og�y
N~�qhmoj�E�ciG��`���~z��q�[��6H��\�M�����w��k���qu_
HN�1����M��ԃN?;���v�߻����oESK��<��1���[o�%�/8d����O��()+W��_w��������E�G��1t�;#YT4[�ؚ[�����WݯRl����
����9dAAq�R��^��Q�K����F�n��a���`������s����%_fth c�����>���iG��N�*�L�w�J��֯_�쎃a����W�a�K@qߗ�r
̹�Y�lU\)�k�Rj*���HX����hZ|j< D �		�,�)?_�:�S,XVNY���0�F�����X�+���',|oɆa(-~�V��-l�m/׊�! �ⴠ�3�s����#"�/aؠ_�QG�_�~�FǨ��>����P\��Y�2?Dp����b� �W�P��������V�Z��$�2��	�2Yɪ��FB�Oars���q��=H&��V�!zu��5bzW7ҹ�[�$��L-�4���1A��hP��6|��0��U�U�wa,�v"u-H�]�.�&	6,�s0�~��G����r�F�	d3`ő�lD:���WT̪1��$�3�K��&5F�/\���q4�D,ӛ��|N�J>WN��B�؆���&�r�HƧ�/���zm}��5Iw�������s����%l�; �Q��0�ùm��zպ�P@gSW~�]誷(�p։G�U���������X����x����Ķ��W`զ�~�X�C{O�L�0^ܶ������~���r�� ^�݀��8;wn�����8�t��g���ٍ��@sϛ�������>�����҅O�B	���Y���m��S��Y�� ���mΙ���5h`0U�p��;]:��F�?�L�V�?u7*eO��#xq]/���w1�,#�/!j����������-��uh��Nr*D0�@0C���#���8C	�k��N}��r�~��({��_�(.�����7�z5���k���q�#��zɘ��cx��'ዟ�4���4+��%}�eL�T"��[G��>u�Z[p�9o�G�}��ct�/���~�3����w�O���H�_��ɇŰFm����P-fR���`��C�'j�Hw������W�ج�j��տ�O@��-�U�C�����s�OĚ�+[ܿ����>�tjL���XD
]�������	P�ݻ�ؿo@�>�]� [Ѱ���B$�c��Y�%E�2Mc|JS+�k�Q���j��T-l��!�so<�������E�t�^�3��К�#�'�ʪ�R�DT��s�N_X\��FW�����	x�ߒ%C��`P��%�<%.7}�&�6I_��q櫘j���M�"hx�q�����v��7|���qBQ�tw"c�\��/�`��)��q'���Q@��j���� ��,ӆ�'��9L��3CJDAT��t���kXs^u׬�"J���arΩs�9}r��~��T�8��Օ߰]\\�}�N����y����e"��' �z4���hB
@-�g��0���z� �?k9n��՘�i�kt����蝹k7#��i'p�I����Z�4,ӕu[�)t����-~�ք�,�%e��n$�ed08^Cˏf��^x&��&z�f�ɐ�f�R�����fj�ب+��aO��g>�ŉ;�{H�#U��8�f]	��*����}5�ă.�|M-a�9��JK�����ٺ��R�B�X�"�v��� �;�ٳc-���]�����ZJ�aE�xё���]�101��0�'������X��y��E'��?���қ�����F`�����n�<G`���ڍ��Ti�ؼ?�Ƿ�a��a�FDf��q�8{y^�
\r�R|�C7cnw�h@�1�mГ}8��0w�"h���e�2��)ݯ �2��_�=�6��3�=�R�p=,]qV�p">��Oc������)5/�=C9�+���Ru�z�R�Li���/i�ˎj�kXޓ��Y{@]��`������p�)m�"��i�J�����8����Â�_�r�W݃#�4m݁A�H�a��8�ԗc��`E3p}'��4�1�o��K/�7>|ӿ����o>�~���[mho�`ْ^|�}������.�Vԣ�=����A��p�	���+.��.;O�S�R�ڂ��==���ߪ~�ۧ`�:�[t���^,MoR���2��jC�E�ť+��aZz`%[��%�L gQ�9D�H�#Ѕ�m-��)?춸hk��Y	�d��xr�qĵj�B�DT�'|,xK�.�)��,䀹�H$cR��-c���*H'$�r�
���Ր�9 & �5a"��]���ҹp�)�&��
�^���
�%�;�v�涤�r 	;+<7�L�0�� �@���_�Z�� �1GP�qP1���&�~[���ESX�U��ږ�Z�)"����_� ��læ�;�+�I��z'��q��f��dG���K�AѾ�,��_����b6�� N�P���-+�DD9�熰pn{�Ux�˰wӓ�Zetvv���_���yn,;���<>�����F!-�njA��U��
m�	�"��Q�w�|#_O��p�	���O3�Z�,�o�h���lVr>���ʵ�m��M�e�5t�v�|n��x�H�����.d�
L����]�zt��h�+rMIq��b2~S�0�$$���Ӭ��t�ON�L��P,Ղ �ZM*t���?���<vF��K�I�l,]|�"�n    IDAT��uk�K~L�V�@o�s�՘�2�Ur8�� �?���y���� ��������X�}���ᆓ��PLB���k�a�&���e�9��-�hq�y�82����R�TɎ>d��cN8���U?tp�r*h�MT�F�н�D�f�IQ�֠�8���+��|w��)t�={G=�Z1��.rU������Ӈ���a<�˯Ao:�Bg{��8�K�x3:�#�hG�BQs]��tc����8v,��l�S��-�w)H�&�F���W>�����h2���s��T�AJJ\�&1��d�(%�P�"������t0��Q+.�����g��m�u�^������ʶ/�_�s/z�	��?��i;v���ų���w�����i88��C��W�R��c��q��RgE`�chKgD_��3��b�J(�!>����x@ݩ�a&(�e�:��o�j@�x5B(�6(:gk��3�ɧ���N<�hh^�z�rI�͓����dT�e9���L,X8;wlA2CK���YBU��Ш��Y�����N��ف�C�Q�LwB��O,�C;���P�\7�J���<��fm˭�HG�	����~!�F �4�K��t��'�Z�JֆRB��>�,����ETn�v���%Bc�_��l��HK�ed_,x9�����ӂ{��\;v[H$;�+v$*�H��<��q�nѕ�y�r�f�6�R��<-��x��I"|��Ak�T����C��z�<�K/8w��jtZY����t�a[1��w�5L��h���>L&Ek#m.�i&�Q�z�ׄF]���*c�%���L�izʒI���2�lx�u&���s!+ڙC'��Բ(���]���_<�M�hD:��(+�*������AM5[0��V��à����\�J�e"i������Z�Q#-Mr�H)��=��T,p���(ҙv´�t�FF�h�kDD��h�04�eK�"k�[-�3����o��o��u�6��O�L5SĚ�83�8p3o���u۷�j�&�������X�c�x|���3�Bi֋��8��98��n,�԰��3[�Z>̘�XG/N<�"�,>�y{Κ��jrt7���oa����4j�t��z��%G/��K���!�mE]u�쥑���u8ʆ�ًL�l�5�p�������ga��i�ry���]���կz���Q�Eo�����*43*�t,�0��Aꑙ�#������_���~�e�st��ޙ+�#:SZ���|�F[g��������.HI��Q�{�ŏ}'$���R:;�;��3��܍z�G������5?�)�����[���nۅL[�5�h �ًw�z-����Q-dіjC�,�k�nʩ���n0߹�ⷽK )�����"�ގގ.����۶c�ӫ����
D͌]	lzI��"@ܴv(���1��/��F)֦��NBS,`�?v.���[P-�����QH�^���o��T{����3���cy&����MHx{�Ta�NM���a��C Bw(.�|E{�鮅��>՚�M6w�7/���C�4���bfB ���C��$��\�'�a�_;\W�q�P}	E�Ѡ0%�笠��k6ZC�Ϗ�p�XB�(0���2��D6;%�r�W�؜��u�L)���&�Yx�*�T'�ši���2�rJ��xtO�Qhd��,�3��c��}8��v���B/�ʃ��f��F$���ҕ,��Ð� (h�����e�g�)���RɆK�a#���j	@�q�eF$���+u�E�9��ք�J��xR�RWp�5��c�𛕻�u�(��L�X��$���7	�U` � 	��q&+iZ��u�6�gj9�S��$ �����!�	����5>ԑ|͔�%eڨ�'���s��ƃ��X~��y}i�v��sa֋x�������o̙���?|����?��wΌ��n�[�Q1���|T�w���mC���p0��3�����#cT��cf�}��	m~
I~)ڐL�d��q�Uh���:�GW+�<~�woA�\���j�}�|+E����/�X���#E��a�Ã����l��.����W�P�0��N9���L����]��Z�$������}+����?��̨������%�Z�DS8��S$���cjS��O��^ئ��PKz{��e�ι�:m��g:�z̀6C�"����:�)���k����Vݔbm]x��?�M�G��Zl��S��g��m����[Q���QD��²Э��X�|!.;�C�e2;��=�������@,��2Pkzҝ��}��jM�;�,FW,����@�.���0��m�HfԀj֨ÅA7+��'�5�|kPإI��$�Q�
ys�r̙ݏ�{��i�Ṏ$���E�njxի.������m���D8;_�"�#����}����.�M��A
�i�:$A�'����'v�v�H h����Գ��C#6��! If��A�'��v���xB ��)���N�#��<CiMP��C��p�0+$즐��Ef�u]��!�̣6C��\	I��(�	e���OB�t[�#u?�F�jObth�Lҙ~�U�G�0�18,��cZH�wH7D���&T3�a�ӌ�Dpm4*0r#��%�����Ced-�����EK�"��T~\r�4�:)˅BFw6ORÚM8�æ�;���Jrn�D����'�(dsr��.S`�l�=���3��g!��/�o��݆	'���;ىj��H"-�8�sB�����J ae*�D<�8����k��$��er�k�/�qwS"��=�Nf�q�Y�t���򚑤8bY�����Y�h1��~�:�_�V�n�ፘ�V�j�{���R�O�m7���ӎ� �ӎ�����F���T�3��+�����c���;��L��2t��Ǽ.g5�.Na�>��]���x����u�.����Y��=gթ�ʩM	%�DSܰ���L)mM�)����A�x�i�XiGGߑ8������fO9��d�����Q^v�]�j|���vd���#:{��ٖ��?~�硯�V$&t���}�)�߼z,���K����Fq�׀_����v�l^Z�08��.�=\��з�T�>�v�D�MR?�^4K0�c������^"Ǳy8�j��w��Ǳ��L�<�JS��{���iM�1:����i��'Ԃ�@|����+z�Z+�k�b��������G�l����W�F(z�&��Դ1n9q���Ը1{� NX����^TA�Ơ$˃���2�z���>4���߄�h�:H+Z�G"��*�;SߑNĥ \~��"(��&�V�*%��r7�r��#�\�O:!(�$���#�o����ػw�[�FܲĒ�֘v�
���<�p	q�:��Sa�x��8�7���	B�4�逿`��5p��.:!�$��O�xRB�UH����-`	u)!����E6������_�����TaG����
�y|b�۬�1uv�`�TB�	4&�T�R�棫�O
�];�bd�.�d�����9?���(� ]�0"��^"��FL�C1��d7�^GR9�&q�+��Eul�¼9�L���gs�j>:u[
0����6(짃s]<��A��6����ف��8^Ip买-�j)��Eb�m�H2����|ܶ0<U�p�Ư�ډy|7�Ѕz�z4#]�߹
�DR ��Q[��'��t<b�.f޴� a���iRAٽ�H����	��a��A�n:�!c�� B	�ׁ�|�<������u��QD�i���%�=���k��Q���=x��Wbv҃V��9/��`��}���_�<o��_�����Uk6�z�e8hAGM��9\�=O����Y tv�u��K���%�8��G7Qڿ(��Z,��v\r�g��g�^ث���4i7�nՓؽy#��;$,�k6ШWIZh�.��&{M�Aj�q��8~��ZT�ʾ	=�����vf��8�c���v\��#�s�VW�{?�>��B���Pl꨺&<� .RV?����s���bU�F����knEz�2T^@�0��2
�mD�&��$n��2��s��P��h��}��X�y7ں�Q��w~��V��e����w���%�6��r���M�;YQ����l]1�pw�"��;�ھ���u�ac��!���>�њ�a��x�&,C��9��.6��F��C��0�i�W�c��G�Y�mi�Z:�����O�U�Dw&�ޮ������N�X���$��y�a<�ԓ8��cE\^��P*L��/���5)tm��8�cD�_��c��>��LLL�S�7oڊ��A�Mfq�NH,�@�R=��`!I-F�M�b<�l��CA��]��Mg��$�D"A�`(:��|=�����*��MSm$T�]�i���Kr�tr:����5vkB���f� ,��u�t&V\���b1R�4)���6��5k�,��$O��
'�v��݋ukV!�y(���W�$��[n��Z�u7�HS�2&r���Z�YB+���� 2����d�`.;�x���sј܂��>�cΞ=��(ҡ�u�~vĂe�r?�)�0w��0���/��r��.�o�R���J0�?���-Ѵ ���k�9��@K9�(��Na�b�W����ډ�ы��e��b���Tf�q��a�{�Y��{�mh��.!�aKb����T"4����y#�f˒�s��Ͼ�v9Jy���a|䓟��T�d���/^��XL4 �Qs��ٸ��7�ì�+��g�t@fʇ��CG��*(�Н̼of�RF`�s�U�V��� �L�`��/�*Z����_�5�����G�`Y��LkJ��a����%l�J������y}�j�=@<��5.6�{k�~�m툐�O^7g�#dB�h@GSE�3�H��;߽3~��z8�N[�&��lP���pj�8���[ߊW��B�5VPZ+���:��/���q�x^-�m�מΫ~�3x��Xt4j~��<�~����e���1_V������˯�]��uYU8�g]����Bԝ��o�o���h��������^w����n@{�|T����+چ�!eKc�Ē�>mo��OaiOF�q�DN�9�J���C2��ʂ6�" �K5��-l90�?����Е�V�Uc��/I� ��&g>�:E���v���b64�G,A9�E�Z�@w�����ὲ~�v5I���!$cq��x���.$�MN�a��uBYaM����P�,Z�'�|"r�Y
S"��z�D�|	7nā�Rh��m"B[�iѸ�#���N$�R=�jv/X�
uk��������NG`�K`�uׂ�Ep�-a�fz�Z8a�!��t�&ȇ�A!
�Yt���tHtO����7SH/
]�x�WL:d��,�c���.Y�ζ����a���҉(Ҷ�ի���{�\�.~��54�x:-�m�4�ȁ"��e,p�b�k�$ٛ�]�����߷W��4��Ɨ�>������X�={6�;�����\�cQ��z���1�z5[���>��zI���S1* �o��b�/q��6"�ތ D��[�Y'F m���DY/�_=�߿o��9([��x��G�J�>�4B]y��Ʒ��^$.q��QG"�;;����:C#f��A�p[u�"xr�B���l��L�4E��ģ+�����u�o��M,�7m��
 1E�u��ٸ��W!�W�*���_�w��q�����Z�����͌�>�`��e�h�� �Gk��o�c�H�Й]�,`A���V���(2�>4�w"���Hc��Hu༫��y}��ٝ�U�A�Dt���Ś�O!e���J�"M�@�UC�Q�oF�	D���^|
�������14��*"BPjt~��'�FЕ�brb^����y*��s��9mϕ$Б����c����kŖ��P-)��>x�<iJS�;۰{����C���Qt��sB�EuE�MD�<�y��xÅ�CU+0*.���ko��k���V"�=������ylDE-�;����Yu��u�{��Z�D��[JU�
+�umg�QGt�k���[G�-�F��1©Ԑ�-����6���T=�+M�u�@]M��JR���u#�&6�����~�?Q>�n���@�M�{�&E���kq�=�`*��g)�)E05�tuu��SO!4-x��X�z�tYX��Ri�j0���P$t!��cv��K�P��e�������@!�`9!\�O���X<���]�p;!5+;�ӲB�8k�������Ҋ4H�:\�C�����L�Zv���Ŝ��Xv�.�������?���z���1U�a���ާw`����D�nEkk��i�A1lѢ�Ƈ�`�Ӆ��@x��F��+�	4 c�ۿq���ȴwu�]�D���
ޕ�*��.���ζx�
Zv+�QX�P1{eZ���	X��t��X04�i�B�SA�$sW8~��0<YŔ���o���
'3SH�3l��lL1&�)�
YD�:~�;��a8E�+.Yt[<�_۰X;��r����e����\ϕN ρ��Τ���R�LFc���D:���y7~�ȓغo�(Uģq̟3]�֬\�#���9������u`4�x������3߹3#03���<<3w��6@�sE�Т�r ��=��S��ුS�їP8mA�\ށ����"Bg�I[�T�\����?��X~l��[��Sw�}�sغa��.����:��3�f�셧�!ڳ_��S�1�BͷPg;���А�@R.�'�P΍A�[8a�2t��G#�%#P䖛��q��/���8�� ����qU�tt���݀\U��EGa��(�l?����y	mC6�l���oG�}@��N�g-i�IA�aBy����o��_q.@�L��J�=�ѪOa寿�����Ώ+ڝ2�����*UM&QoV�1���"�B��D�TEg�Cf�O9f)N;�]��Z�٦ݷ{B��=�pE�kǑ���2M~*�U2sK{PЦy�\�gwcplH�bL/pB[�X\�q��t�����.M���Pn߼I�ܳ?��O122�����޹K�NG��fÃCصk&''Y�*e�B��"B���+BbD�ݑZ�#�B�b7�`t6����{�Ů � �<��.,�C��.����tQ�f��iSA�_�PP` d4!�	]���a�!Ha�"t�
�(a�EtH�
חk@m�4����JP�c'���.OС	���-����X��װh�LLN��;���/���YB{�?�]�8�g;�<�(�,�����#��0�0�EH4� �N��x�U���4$WF�\XJIG��;���<w�|���ݻ�x]==`]�����;�l��U.�Z�K�:;^�dLB.)��y�@����F�z���-�V�]�˩���D���X04Q�h3���v~��6�틑��h��ݰS$�JC[[�3Gv�_�N;z���j!���|�{ulضC�
GF��K�}"# *J�j�)�������ZMlC���������c�Ȕ$��:�Qk��YQ,���LV?�l����݆�����4��^z��GK��������<����@ό�_�<��ZUm�i�<s�F;����G7b�X7"�ʸ�З�q����~$;P8�	݁铳mC�Rx�5�@K?_R�����"Ќ�
��x��o B]g���v�N��mh�I���b�9RpD��1ہE>iD�:�dn��i�D�S�۬ �4��Ī(]
]�f��3���&���?z]���κ�J�Z��_��\n)�����=�֘P\����'pՍ�F�}�������(�b�1 ��y���,D]jB�M�V�A��LM�3��"�Z�4[
F����*�Tu�A��� K�ut�KUt�3�IEq��NǇ�~ɡ��{��S�|���[p#)�̚��1�u'0�e�8+�a-y�I�Z0Ϯ~V�FjJĵ����W*0�d    IDAT-�ۀ٬���ރ����6xp����xꩧ���at|evZ)����j_�g�V�,�	���s(�E#-�I��%H	
�8�΢�v�]]=B����*�4��%(���,RÎEX��|?;
��0�$�b���$:� ���V����APH�
��Q��B�3��b�P�vjD�<mҚ��C :aq.B;j6���NA	_������Ӄ�N:	�dL�:S�ʍ@�H�ʵ�s��F�&�7{�����(zQ�tcc�J�:�h:C���<x�E�Cs�#�ʸ�:y 7^u��B��E��$m]�=�' ������nL٩)�zD�(��:`3��wĝ��h��IӔ{F�3)u|��5��g0��J�ء�9��Kw͠����1P�~abl��ᚍ޿�xdZ�y(iq8f$ ���h"� �q,�y��|�榷`Ao'�V�FC�e<W����=�*�t{�5'�D�˥`���YA�G�h@�mZ����@��M(55hVD��%�=��s+�
�������w^���U��+_x�L���%?s�6#0����\���s��k6�:)H�&)����l�<��eQ�"Z��B����E�����"�؆��琱ZHEMD�JM���& ���㧠s�&G�+�_Y��D��c�
���-E�TE����c�,c'�ϫ��(J��<��~$�� ����l8�e:P/׃�UJ�":l���#n��rq���j�H��v4"bͥ�zq�uW��3�h[�Z���㓟��Om�k��G�Wx�_�Ysum�hC��v�5q��oC�c6���Yx��ʬ��Qe�x�kq��^�Z��h�����[>�Y��Y�Pʏ`����F���tpTg��y�kT�e"���	�����D�� 
C�������{�u��?�l+��G�����hN��o�V��cM�p��g"[��歛DԪ�ę�������Pk�j��Ob�#�!�j�L�Q�B�V���A)N���g�1�u���* e�N��A��A�o��mli��b��5�AXtr���.Y����ƀ� H^�t.����vB[\z�qH�4�C .�~�n��<H�i��+a`��]�P��u��� �C���;6��1��vSB�_n+|o��� &�s�#σ����5�+��L�g�}z�{��0U�F����p �NF�z]�:����~���]���1`�14yihRwK c>��&3-|��@�0��|���\���A�,���H���(Ml�ٕ���k��B�]._�=-�C��(��e�� � �{$	���8C��HAu\��A�J��B�Թnp�L�W9>�e��8~p�Z�����P�"p��hS��B*;AM�S�@[<������q�K�@;s[��,�z�֬���-L����D�E a��q�ZС�x�<7G��]�tH�HM����b�+�K���3�ª����Ew{z��0'��+M���$��9|o��_�� ����6s���<�j��,�2ZҮ�2~t�Jl*v��#�`�8�Em	\v�1��7#�#�U՜�sߎ�e�\-��4����_�4������֗�5(��J�׳��b��l;0��G]%Q�G02��H�	_�zA�&yI!A*�
P#hr0�T��p�y$�f�鐮�l�LO�=�(֘#��"��^�ܶ(��+q�K����<u�COࣟ�6�x��f��d�^���{�X�2�q��*���]p�T�.�S���V�B�����߇�N����$�f+���n����w�z ~�N��5��
VD5mWaR�[�ޥ�z�U��'$������� _]��L��BD�Hj-����K�]��o�T�m��d���'0R6P�Km�cq��#����A"�ma";.�.vqP��d�3:8��9��A5�����^�ꗢ'a�Z�@g:����
y���E�X�v=V>�4�9cO�社����۱}��C��03#����d�]p3(�	,��)K|_@��0��R	�Y���,W����S�ف���t����R�6D:,��&bwz���!���Ӑ"2��HA�����c��T���}���'�`q�����q�B�r�'ʸ�C�)?s�,b��������1{"&�&wsiT�38���R4���.]V��b�nE����Bid`���V�JN��|�c,�݉��p�egᖷ����&�F���G���3A�������9wG�.ߎ�ެ�!�@�`��%tt)�H��R-ǕLj=b���q2�q�<��Fv���4�bMC����~�~�jN|�t�~�l8P��i:|�D�q�#��ݵ]��z���^�3_x"��cH$"&j-������$��`"_�l��E?�H���, �%R�,F�	η��5�<����VoW7�����]{��1?��e����k_�9Ini�8}&��y�*���_�� ���<sz����?�F&ǥh�>������a��q8v;L&��8�EI��,m��(�BR��]��s���<�W+� ��� ���JS-dH�����_B�R(�r�=��A�l;0�}U�\��pp���rPJ��o]~r�L�}�x���3��<pz�I�2�����eK���4������Y�{�Q����b�^T���~�����h'��	۫�럼	o|�<mK�QC�ց��=��Y�(�eqL�;A�kh%�3C$�O�]x�Gi�U���i��Y��3���ݨ�'�ܽ��4*����S�O��_��'`��� ���W��އ�$)i�.y��ۮ@4P7�^����'�mF�x)/���d�PU*5vRt�E(��J�A#~2G��`z6-���f���ťM�����^�Rdڒ��� Z@��P�V���D'�nZ,v���H`�Q+��Nd*�?�[� �I��*�CרP<���Y�T�%�K�I������F�� ����8��u	$���.��z��`���6���>:*�%o n��s]��C(,�Tlۆ	4�q�k��)�����oaaH��p]I����$���s�}ѢEؽ{���B�_�#é����}"��Ԫ@���43���4��4�M�|F�#ψ��I���8�Sf lSr4�zqSGO:��x����;���׼�\s6Fv� �g�gV"�M�ʧ��z��zD@?�$��UNS���dt.@��!	D��fE��t��3�g�L�Ɋׅ�P.t��d�A�����(~�r^z #&T�V�9$�K�oѵ�|����-�4�+.� �����E��d��߫��:�e\
-����kAF����J6���:5 	�L�H�|�RF=�-�FO/�z��k��%��,_4�]�:d|��Q�{���J�o���gF`ff ��=03����m;�ä�8��ף8���'����h�4=%_���(�#��K{�%I�彈�cH�X>9�����/���F�K ��ゐ��s*jBx�;6<���B��Q)�r�h�*�8�m`�n���0UְsN
pN7��Ɣ��B��e����9/;_�܇��[�~�iP��MoA���,={:f�B��1>�E�-#������|-�=u1�Z
x�?��<����h�ت�_|�ﰠ��b����ͣ���c֢c0��B���rA��LO��'a�&�S�{˵����ݥ�G$݃���lٗ���\�懿�V�$����Ǖ��ѧ��YG#[ׂP���7�5�=@JMIvF��q٫^�����X���M{�;?�	����끸��"�M�@s�%��E�	��
�,2YM�n�#j�k��0N8�8\��s0��O<�z�Q)�J��h5hg�pI��ڃY}"8��|";)��,�ŉ�:���n�� ����sI�h��>�[��y�a��E�z��¡愀���@p�!͉�õ\/�g��-������᱅NKE+XB�T>�u���D���!��i�P<Ҧןn���C08ri����?�/"fߗ��n_��P(�1�ƥ%3]�<�ju�Q7	�<Q��|4}p5�������P�]S;L3�e�rԋ4:h!A
T�
�U���u��u/ƻox%�w<�Znɨ- $�L��k��bH_Ĉ�p��#��͖L5�|���M"v@����Lw �/��0؏�#W��j�&B�:�5	�M��h�?��1���~ U3!ᤪI @0D��g)��&��}o:@�T�qKᴓV��7^�7�t�*u��t�;��"i	<��:�(-
����~�bw�r�,pc�6�|�%�>��f���۷�D�N�V,�ǭ׾�STig�:��) fF�� �����*G`���4
��AZ�2"؟����~
��BUK���L�Q�+�sRx�)��r;Ю�@		�H괕�㌗����K���?�3W-�Q�F��2�)����;��Y�mv����X�v���PAR��sU���UE�@ʇ��ǴÑ/����.��B����:�O|�.��_<�m�G�5g>bm�ˌN���V��]7^�k/;K5M{l�����«_w=�T��u��KU���-���&4�O�Wo���Hu��x(V�"NmkK�Z+Bc�ů��������6���cl%�e�p��>���9����"���K�J,�:���^���B4�$<�>LvT��0G/S�a����/:�|��ږRKœ�lĭw|SZ4%4��6U0�mKA�@�,M���7lJe�B�	(*���&lUǊ#��ַ_�T��]?�	�[��̼R(K���*4�uD�'�$���H�Z�On�'�#3#���G,x-;�#a��'���A�x((���	�v0��dr
�CK^�a6Hh�"��s�B/�u���:��°A��LS�'�@`vExl,�C���@��|�1��Zt�
��mp��~���M"��;&�f�� �u(<?�;�9t��߸�\���!z�2�Â�1+C�#�L����g�˛�R`�3�,�uxԂ��r/iv0�SN��@SYyrc��D
c�qÕ/��q	�=�F~
q[ �̤�=��!��I-������߇��^̞? ��f��H$p��\���V�
�%}��*f��uq<���K26�F��X&�QE�Z�ZW[;J�j���(~��>��y��:�H
ʡ�V@�#������#a&�\�Z��O���L�V��"^��(m�K_�r5Z,-�jp�y�P!���i0�$Nwo�0A7%!~ά�����ƍ��h)8�
�Z2���H��kY����(���_�3'53���<<3���6+�oR�$��l�
�ö�)���&<�y?jz
-_G̶$@Nw��\rƱhײH�1�k%ĝ��_6y$�<�����8_X���JW$�RP��݇��-,�E[`V�L�J�g6#��?֍���R+�]��(U���&�  �X�H��F	��x%���7i��+�Ʈ��־��G��~v7���2mؖ	�E����ȃ?F�ʅ*������}��ʵI��Vs`�*���mx��󵭹�2������8�Ξ~)F�Mg���f� �;�ٿ�t$���E���z�o=�M}���X�	�ɠ��7��9hU�2���3��:鵪dv@K�H7��H�i�w�f
�3`z���鲗�淞�f`���W��<�Z��w^�6,x4�7�==�D�%sfa˓��+�a��z&���P�*�	7�p521O=� 6�_#����,�
Ų�R� �������8�c�s�^L��a/"l��E�V�0�h�w���qVx�RW,o�@�d~nU|=ԅ�T'�E8;fa28���H�r�C9!��@H�
�sj��*�ʇ�T! 	�$�ݙN6�*a�9�ǅ !�R����rſ�`�w��q��B�c��%Ԛ���Kܠ������dj�^n�ך;bҸ�iٰ�� ���R<-
O�ॡO���[hp�?��g[����B��9(L�CkT3t��%��GPۋw\�
��拱o��O�1���]�t�CXh���g:��=���A,>b	z��	��"u�I�NK(��R�z�|A���-K�ڤ�G�|�\:�$/���p��B��"W�B*�@og'�F���W�~��~x�$ �N�y"l�@$�J&Gb0ЛI�)塹���;�I��|f"=҆�.��N��j��갦)s�(l�ր ��u'�9si[tZ���ޅ�ϭE��������W]��Hf}
�>#B�) fF�� �����*G�gWK�߃�׭8V�8�U�'����i0����D%���ÒvW_|&��rrH�U��QK(=��Ypw�ؒ?���N�RJ5dfݶ|���R��H�+�
l���4�m`��QԑB�eCE:QWqlز�"��|zI���4vC���<Sn������j\����k��Qu��~mKQ�\U��SC�dR��$qq�r}�mزk�?�,�� �1��fÎ�a4���͗�B��EU(Vp��هƇ���%_jOS�EM[s`L�.Eւ��}���m� V�W\u���i.���gqr���*)E����
^f6�VJ���M% ��{7�h
�Ƀ8��G�S{����_>�o��]����<�9�,��&;�An�ec�X��?Tj�ƓP�";'��hl��Z�JG,쇍ʕ<��Rm���%RR�;����K�X.i۵z����m��X$*3�����"ۢ�Ʋ��zM�Ti��U�3ڡ����AHl$�bU��0:.�K�Q�fpp���6�0����B�Ц�{P�'�/�ɹ}v����b��C�A����mR�vJ:C;��89kO��c�k;$�Υ.�.�np[BiA�vb���֭�j�RI�Qd2	�%-����h@�mi�cp�.��.�kR��-%l��aC�,8� �@���t�JYhQ�qv�e�얱(�\D�&�c�x���=on]�z.���7���4��.vi)�f���DV�����2�@\��Lۀ�0�R	Q�}ݐs�M�$���i�.F)����dp�}%�N�����w1;&`�Ҭ"��3�F��Ɨ� �[=
�m.��~e%�T��G�S���wS��sv�g�כ@���/-.��B$�tDc�$<=�;|7����b�AZ[}:A��<�l#�OR�4αLwA�9ؙ���u�u5�¢���%�j�j�FDdh��y�+��I��s^���U~�Μ���#0����5��_�<�n��5��q��k @����{v3J>�8�j�����B�����Fu��A��EX�"�21�2�t̝�Sλ��C����^��K���2��ٻ&�}�~طWhC,��-�5[��S��&�����D���|ӆo�c��`�$:�P-M�S��}��24$qw��������{�`��c��`#��	-
U��pk��xR�I��6�����_��߻-=�t�|���#ڞF�+�+�o<e��qtB�w.bXMÊ�>m��(�ہCQÓ��]	m�h^٦&V��Sm]A���Q|��~��Ֆ'j�����;�L�5��o��G	%��mI-��$DШi��@:�Dap�\ч��Ç�`���[����ޅ_�}?�ݏX�T'ȹ��*t���~��BL��[8q�2���>����8a�mK�
�xu$":.<�|���pԲm��A����/v�M���ի���b׎mHD#�?o!�^~�GPn�pppP�d�	6�������eaMj���:��K2mWҗ���xG@�9,t0t�
u��gA�a�F���{8�?E�>��N�!x�����ì�i�8��b�
9��p�]�����@���ҙ�A��s�CM�g�s�Ν;u;:::p��'K�c�R�6m����	4[u,]�g�u�hq�t�����T��Lg7��;�g�nlZ�V���Cӥ������tC�5Iϙ�X{�''`�&�Fh5��d�c����<z ��"���cd�*4� �Ճx�     IDAT:.v\t�v�q�
Md�Sr.��M��$��U��Ȝj{�8N�G�R�7�I�c��E��NaxdL>'�IZ8� �|�,�Q�uv�x��X<�t"G�a܉�?�Ol�������÷�݈O�a�U��Tu~��c�\�[n���z��I��9\�<�0����3��oC�._��r�\�
� q�
���=���G�"Pg�;�P8b�"$��|�q�K&"8�����^�Vn�j��}���9���-:s�3#������7N3k�/�U���_���oD�u0�U�����m(zq�}�4).u߅Ѫ"Ҭ��OòF� ��0��"Rz��p�2ݽ�����[;�.ņ�Z�_>���N�]����o}qN��? V��H�fS��aG1��`��1�h����X ��`$[�X��B��]��}�~�x9M���=w�wJx�K^�w��v,�E��h�R�z{�(�����021��W,ж��Z�~�y�O�v�A�v8t�1L�{�*�x�����o~ؚ�=WP�FE,@���,��I�7��Kۗ-�f˓�aiOZ[38��ٸ�<�4�mB�3����m5�C��n��#���v���x྇Puu�i=l&$ڎ�p��P,�X��0��>��y|㫟������O��a'�I4C��?���D�Ϊ݌vt��,����ݿ+^+��Yf]f���<$M�֛�Ň�u�z?|�3�S�{�Oe�x�b�F��Cxn�Z�	��)mve�8�b�v |KGoo/&'&��bq���8�l۶E
�J�?66"�
���>Zl�x�)�`���$P(�X��Aꨣ����ر�P�8�����`lڴA���:�b���u������ sE���r��q��u�V�?�}饗��;�̙g�)��<��#�{�W�����s�x|򓟔O:�~�%� �뮻d}}}r�,�	Tp�\8��u��ͷ������J�P���3�N�v�fDP�{��bF��7NɽR�m�7LX�mp�)5:�F����5;���?����2\��ax�j4����f�� �L�$�HD�����a9vm�(R):np5�gh�۪�e�x��/�ۺ���+F�0�+`���H�S8樣�ު�j�T�k�5=�hQ����$-�aa�b�wދ����'{Q����)�QV��"���`�R/����7���*�D�3��ޚK%�J�%[�l��<�`�������@���/I�1��ˣ��W 	cLc���A��Y���P%�j��g�������=� �{�ҒTu�9��3����7���;PH�L錅�|�s��W����L	M��!]�Ҳ#.W��P$Yd�s.ց�HM�S0�Y��eG������g�AO��g�y��\�em�y��x�ݷ9ۭ�Ww\�~AJ��a�;���o�����&;3�3;/��#j8�|y�\���}e|w�Ql�q�V��]�Ի" ��&�_5��V�`8 ۚ�^�`ڃ֞���L<�r9���04���`�0y���I���n��/Y��s���,t�����4��Ɖ�c�7�� B�� �m��>N̵p�T3Ma��Ս�ccr����&��f�w�
��Yj4��m��6P��A�ހ�y�����/�7V�X��n�^����q^A�'G[Q�����ǟƶ��861�4 ��I����H��М9�p�>������lF�ꬦ�8њRj��t�܊���������?l��ݗæ-{ #;_�/W9iYJ��&��jT�І��1D��ƙ(l�(�X��D	=����ܵk�}�
��=����bdRR�p%�u�,�tAwު����3<�����$Y������y�{����/�C%��r�>���z5�����ƞR���w�^��oF��b|�܀B���*�B�8��d�͂�E>�+vX$�u���^��_{��RLn~��XīI7��o���o~7�|���dp�H�a� �E<��W`��R�n޼Y��,�_=r��}n��׮;���133#�-��"��{��q���a�er�	�I�<���h^�������繿u��I^
��E5��Wb�ƍ��Y�v-��y)R	z*J>�������g9W���Q��+<���?�p΂�h��/��ū{�Rkcz��#c�hr�Z�C v���|�`��	v^s9h��Y
t�w%�Ў���h�������=�11���I2)���|��u�Y��5P��c����� J x�P����R�sS����i[h�-�9� iUL@٢#�i�=p��1hԄ�,��9�w1��p����?�u�p�'�u-���Rߨ����rj��Ԡ<�+.����.��P�TE�N��2������3�H���#�MD�;Ie(�Z4�l^��V�F�i��G03d{�Qi9�� z��O.<w�K=x��g$#$ej�z�Z��[��rZso���N�3�m����tn���3��Ot��N B�>�q}#��{����Ć��4�x\�#�8�tb�E$�.�*�_ه�.Z��?gb?�:��RA�|�B��~d����0�d�|7�G�G:���Qəq�-p4_:-.�t�'qrlS���׫��3�y�qF
85���T��!<��(�f1]v1u��v��[�>4-�.+�z�"Ֆ��#�G:�CO��r�P�̈�օ���^3����P��zhq�������Gy����hy 2y�{I([ļӂeXpk�( ���ߋ��]��~�ā�'��UBWW�T�X��a�	�r�)�p����xn�� f� �������{c�ڛ�B��S��1��
iK4/��rju�\���J�"���A�@�G�Dz-L�B��U���F����Q�H�v�r����x�nU�h��׌��|��n��r�z��X6܏;n��>���o���9�c�ʳ0;=��{^ǡ�ػ�_��Bx�f
v7�9"���n���_yDV�i�K`r�M7H��Сx�������	�#IȢa� h!H��ˤ�g�E�L11�,1m颋.¥�^.�SO=%c�p�Ux�O�箾�j)��~�i2����p��Yg���-[��	�"=������{�B��c'��vs �/]�T�R[�n�����on�ox����|�3�wBS����x�\���w�[���u����۶mFen{_=� )�;x�f�h{�5��TV:��I�z$�<"�B�.�s�+ bu��1��� 9yx+�i�
Y���*�=)E��0@:�CP��;&������ʂ��UB]-ĩ�I�`�!,�F�T��늿#��yq[� ;���Ǵ�9As~�����#�2Qu"�j�����<���/F��&�[i�C��G!e��[-�i�/?�j�%��58d���Gz�3�^���4�4��JcM�/�V3��m4�JL��JJ�
.�ן�<f*M [���F���.BWW/�|j���Rww��+��{nE�Մ֜��o����O�K�����Fg�@^�'�3����]RpX0	}����s/S��g���~��1.)"����bq�����A��>�
򡇬���v�jk(uѳ�O(CI�kL�1�Aٖ�,8L]�rj#B�	� �:L6�>;'+������|[CS���K�#��s-����W���C��}:�x"�@n��ϣ�wV:��jKG$��,�)���{�m�JS,+ە:���x���m`C�m�J]���℥,nHW����vD9A�E�Z�cU,m�F�#)�,�X�ѝ3��T�-"_��q���mb�J�)��H:��Ta���r
J~ϋ�C�B��t��%�!]���H����!t:Q<b�Y��j3ӓҩ�����ۏ�<�ƥ3�G�|d�������~�g-��W]�=��SW�Y�P�8qB����)�산�bV-�������p���<�+��+��"���.�T CWw����Yyύ7^/] �ᢋ/P��/ʪ��W\-��g�5x��_/�������&�>��P�KS�,EP����֮=[��K[6K��.�:����8���J~��X��<�r���P�x|�w�Gr��|�t�MR\�_�m��&�G}T�-����J�����m۶ɾ�^"�vn>�UI��.�F�1.�/����_�N��u�;p��Ʀ��k{:��I�-0��I��O W��s 	���2$�⚶�A^}����{��ѽϡ2;��b}��r~�����k�`:����>|s7�4��,8A)#
[�M5��&��=L�AN/�d�MQ?�#Ec�$X�q�n7Q�7a�t��5Wä[ć��xᰃ�8,�ޗ�K�"E�"��x�]x���
#t������ڲ��k<S�� �s*H���NY���I &;I�X���x�6��^܋���Obǡ�h� )��e�C%B/�⥗wHgyQ_/V���7�*N�Zc�#B����l�d: ��Dw󇛁���Z��Ж���Y�8r
O�ŶC�pB�{Q�KrxʰЬ7���^z؂��	뚋��߮�lL ,O���Xڟ��1��G6g�.�������*WF�@8Ut��g~1;�XX�D�	ݨ�Bqә�{���!�h�~̵��o���)yO@>G�/`[�\u���
6�+��ct.B��a�OL�UoCKg�sa�m���L4[U�r��,J�YƱcc�����n*�}P̋H3�9��'b����n3�0�A��$�0G��z|�U��md�Y�͖�Xъ��Jm��ʩXQi�-�h|�m}��@V�%y᧯�V�`OQR�:%�[!���9�T�O\H�S���\d�-Z�֤P;��U���'%�!�s7�E�HɊ�#��8g�0>�@�
aj!�-�ʢ�9�U��
��쌀�R�[ A�؉q�Ld���ju�E�K.a7iX7�x� �u�+?{����-wK���\_r!�9�|�k_ZϢ��"��gXx���B�T&��R��l�q�}�attT�iU�a�=��r����η�X�&aɒ%R�W+u9v
��ĩ��1�;6|%!�6l�t�wJ��c'��/�M`�~�z�p�����O�<p��q<쎰{�
�E ������fx�b�v�-X�r)��݉}����уR��Z4qj:ݞ���~�6<.dXYY��7M}�}h�`2��`� �s�vqE��B�~ y8A�>�_߃_��J��4�N������>K%Y���!�G��r�R�</l�a딑5*�RZ���5��g0��B��H�9m�	�	.y�]Œ��*W�(?%�:;�R�uS�siS�l��x=���x�P�Z���cL���q��G1�F��8.�l���>;��0�t�|��͗瀞-���<S����C �/�\ۢ�. �tÒ1R�����;������Ah��lA�u*�V��@�؋�;���m/Ě�~��ۑq�`����.��P?�Wk�]���žΜtf�3�g� �Ҩ)� +���a�����8M�Pi��|�L��ԓ�`j	2�n�}�H�r�����u��j��75��2�e�)��@�ȕU<v7�!���\Yg�E{Hx�M����@t��Z
�N�a���81ۂ�텖��1]uq��$\������`�i�J�}���B�d3X�T���0�\��LCcR4��)�dzFG{K���-_V=��3�������]��J�R�kM�}��La[��-�zE��,U銤ljYԋ�v��Z�?&Dj� Ҧ-@��#��gA%�bt~
UJ9;!��Ez������ݝ��Ӈ$09g��I�}d�y�-hU3'd:8]��P��,��, C�T���ex�����>
�#f���eD@�f������p�e�i�G�D'��sOiX`�I�Et�2�J������U��(V!|@��24����4�D`�� ��Ko�G~�b����$+�w�y;{�1~��W�\�ǿ��z�B�!J
9]ǵ�^+�&X�vX�$�tPz��,E>�P{�&m��6H��}�g�Ŷ�B�b���	��w�Ą ���%��x�'NYAη��-�^�Zޗ��zz�'��Y��E�����m�ڵK~N
Ǳi�&E����c��Il^k��������o���WD��Ux�����l�)�J�Po:���Mu��E Sr(�� ����w��S����:�<����_��߲v<��ܴ ���^�g��@pC_B'��j�Ut�������n C7��'��E3SL>"�Jb��s,�Uke��z���6/#���@ք����Ȥ�Ƒ��?{��|�) �v�^lx��^:M(tTg�0�Ӆ�~���B~�ˤ;_(�y*�鲒����5e�!qPS	��:�9<DV��o��������!v83[@��2���c��s����v��)׬_����f��i��<�tͥ �) :3�#�@���'���xq�����eJs�c�c�ζ��?QE�g��\�Tn4\U���^��XZ �2�\&�[�|��$���aKJ��ݭ"���DA�m�B{��#C�m�P,J!�/v��Й*�)+���I?:xl�-�6�Ps�"aׂ�g1~js�U���D`��kբ&B�[i>�#���ۏ�Z3�&�l�X��L�\�d³�vt�<[V��3�C@��2��D�ym%����h���(~}sj�MX�L��@�Xl�O����D$���O#E��@���9��\r߅*E�*��P��U}�s����ǧCP�Fu��%�Ձ��Y�q,�c|����2�//nh,p<t	r�m��A�{ �{�F���8ni_�TF� F�F{�8��6�s�󹌬�����]$�4��ڱS��F�������XӺ�3����5 t�"Hx���,+��|w�Гff�d?��_,:�$��:]}�o�(� &q�b�?#�P�4(�
���J�L ��ȳ�>+E+	��cc!�ݍO�X$�a���h���E��gϫRP��]��L%�$ŝ�:t�8����kd<�׿�u���h&�*�� P�c;4��;��9��~���A�4h�3�I��f'�e��zz
0t����MI�n)��t-7@S�������t�a�k�B��LJ�y�Ӎ- b��|DHEx���ć�}1��( ����@��AI���P���06z˖.�tr��f�d�G�V��y�a��T�큝MK��j��ʵ2V�Y%�(�W�Y-�*��8g�]v��Clr�����>����p3Ch1��`���tA�`S:�L����� ���7c�@?��J]�LM#_$�Ԃi)@!c&�����,�g(;��}����R���k��o`��D��'F����V,_�bW^xi�,���k7��w�퍈�#���:.X?��@�~3� ?�Y���53[^y5b����r��E�s|o܁m�N�G	>��[�]��D��vS	��f�HQ�6�tQ����?��1�TTE�r��"d���ʟF*�,����N��|�(be7�P��Pi�G�pՉtLUZh:ھIO_ ՍrK���*f�-4��@��J�S�-m�):Wabfw/Y���٦�j2�5/]�R�L�D`��F_s�_І?�IW������H�:ĕG���Na��<mM%a�R,�"��&�LF+Ɣ
�Ό���հ��2���>C�ى="L���h��!A'�ʰ�?� FR�$E�K~GZ�p���N�+j<nJ�C=��I�!an����a��M�ð�4�z[&�X�sa��6�N�S
V�1/����HHS@���B>ߥ0�E����Y\���w<e���IobQH*�Y<�q��R�>�ط��X�R��U���)9_���6��쒰pO�:Y��#͉��.�tN?� ���(����8�Ç���c��	x-p;�75&<w��������}���&��uHZ��wߍ�~X@���+B�Ck_��4-��$9��#���bv�����̏�Z�Θ`H�Ln[������g�� OM໪�@��Z�9��    IDAT��T�$���i�j hR�Sä؆�(��<4ۆ�o �@Z�������qx�&��3(�3�I@���H����hW�ص��9�lt�E��y�&�m+���4^K�'�z�KPS�a��A�j�y�w�:��X&�C�qč�t(�U�s�< �OW>�����>>�����I�W ���)]�8~���Y��ٔ��֞#��b� i��X�eDK%FA a�mו�`��D&_��h4�@�дL����50693SD��H���)8�֮Y�l�[^�.�W��X������.�2�����+:I诙/��@�f�@~�NIg@?�xq����a�A��T��_=�yv^/��ņ�+�R�R��`�����f�jS�������|���X=RD)�A*Hk�vF�bE��ޡ�%C��N';n��]'�*�Œ��&�l	��@�g��4�{�̷�xl��ӝ�"��g�f�D�����]����G�؍�������#��CCH)zq;�*�1I�j)��Q��S8O��V�	lt�KDA2�t��h[�>J��[�N���,*��n�zvKrB��Q�ZR�� @M��()�H�o�\�UR[��G0!��bS����E��f��p�3�v.���S$�0Z7�YR<�z��|6�ma��!�ٴh6`e��Ύ�z�L���X�|1��0?=���,�
�^K�.��QZ��b���,oM��=q���!�If ���b�z���)o��f)�{��R��bĎ����}�s��͕}v4X���D{^��&��v7X�S�΂�ūJL�a���kA �п|8nv^�'�
��@�/#iP�w�,vw�~EV����W%BqvT�9;E�<6v1�xy�x��mo�i`��bn����,��1��q�ԀPC�X�&Y'<�/��r?�K�mD�!z�.�4t�}��"m��B��J:M'�Nm��������B�S��4�(�f���x"��c�E�4�k���>��_�=�������Ө�TP ����Bq�jQw�LVqh��^�==}r�:5���o@��`���P+�q��qV#0]q�
�G��[:����?�/sGa���N��bzv���ŋ�T̢Xxe��?����X���݇fd���汙\� `Ӆ��kI�.]��3.��</ҩ�D��uyx�A$����w}�0D.VH����A�{��Heu�k�Π�1�!j�tѠ,]��b�n��P���W�w����
Ra7]� ?���ξ_�3� ������y^=z$:zbL}�ҝ���[��]G����0��.O쒰���H��6И�-��(��S8�\�&�jQ�T��.ZȚ.R~&�na��<�.�3i)4IY�ٽ�LX�\_� �6;	�[Bͪ��&f��]
�	�N[�2��� ����tu#�ݍl�$V��g�)8׀6��\���elI+eL! ��=w�� )N��g���S�`*ŷp2�� �I�"لĚ2<c�d&%<LWX�5��
;b�I���:,2$|Lu=����v�NG�~.�b�d&��8m;�f�Ip�s�����E:S�T��T�lV(��'�:�$I g�ı�X�r;7~��)@(��"97����E���KG���8vx/,=D>����F�C�؅z�*`�V�J�LP���R('�vNX�[�)�2��e˖��6   9th4N"V�X! ����i,���\Q�M-�8�"~'P���+��q�Ԕ �؍�g8�a��#��ؓ��R��H#pZ�b�tZXs�����on����}�нz��z�'Ҵ�ݐ�wǑ�'���u0��9���E��㡝1��_|��2�)�%ִ�-�&HS�-� ����5&��V�,�_:A��n;Ȥ����=)��}��{��!�
v@x}f���i���.x�0<O%��.֫@o��'>�^���aLݎVk�t
��Ho;�ق���ܿ�0^޼�^|���J��#�F1q�$~�oCw_�h�x����q��~�b##�ܦ�&�g�26}�*I>������?>&�Ij��#�7Un��M|�_�h9'3���Tf�%�]u�B��K��t��u�ivFؙ�t>}�A:e	��y�ߍv[�m~��x��\yH���2
��aҘ	��T-�٦�008���2y�޵G=��[���D�+�`���;5ԏ�;���_���<�8�s�?�<1>�l7)
u5[����/ �%�B0��_�F��&�F���t�L��Gh�i�(l��ߝFut��=Ϣۃ����lHͰ�ju��IP���y�tB�5WhY�z��#"i��R�M����>�&��z1��>X�,Z��z�-4�E�R��;��@\X����ZZ?�AJ�!�$�ؕ�-n�u��x���!�!�Q
Ȫ'9�Ԃ�&"_\V\rv1,��+jx0,,�7Γ!&[qG� $�}�t,(�� X8�:#����3����5��2B_��S�@�-��p��4�xt�qE"�-�%�e1wΪ�y�9D��3)Z�K�bxq��j=.:�,������Ø�:�BQ�mtq�E�I�űy�t-X Sh���^)��;��8;Ԑ�*�2r\�g��.�U�R�(M�B�rZ�=YY�E��PHiZ�j� ����p[�<qn	��'�C�ւ��s�X���zg��F@@p����:ED�$"g�%U���P�]	��@�%�q�
7�N��ϓ
���$c�>F������9&�h��m������٨��+�'���Md���"�89%��,��T�z(���S:mh�O�;���[(�5!�:m���A��U`4'�ɏ�w\3���^��5�I�X2D!�W(B�3�����=�'ۂ��{3R�4̴�f�&���}��H�ݿJu^��ў�n�vʔ�v�-�[u�]Z �r>x3�]��>�O�R7z�%�u|����-����g�K���΅�tF�A��"��� f@��{I�QTG�]O+���z0��%]�e4�,uE��ՋZ�-��+6sF|1	<i�K+�"7 ��:���FO�rZc�������ݰ�YL�]zQ���!�W;o�������ӹ.:3p���8!�K���k8Q�؋����#���&#.'re���\�' 	��'�K��PU�F>i>���JY��>�D�V��R�4�U��*�	͚��ȗ��٨Tk�"^m�Ш�e����MWDjS\m��ʕ>�*��_�\����bz�A��|�
�=mO)Ty��Q�$��)���.�W�	{2�k5'�X�8�ч4��0=�]Z�j�Oȉ��r�/}f��5���hb��$s�X����%�/;),^�o��R,BIP�G70���P��X��"��ް�<�G/?�l�qЬ����!�ߊ�~ &LS�r�ʥ���fD��J��D�}A�	;ca�'���A�x˳'�-����+w�HC�\�/��YTq�~Ŋ�R����⛁�,�%�<�T����,�Yȳ��pE���΁X��N`[�\�����$�$ȑ ��9��x�v/���F0�s�m':�}�*U\���j����ɋ�����I����g�����q���t�22gn�s��&�@��}�3±�s�.������$�F4�#�����u�+���6v�܊��~��V嚃���Ё�9��>��{�]Dۃ�� @x
]�ע,d����l��u����mW-Ɖ��%���:�����JKFP����^|��gp�6�-м�]�6V,[*���;���1��<)i�ݽ=������F�V.D4[�E�)��|qs�"�\^:��f'f�8<��0Υ�2{�P�%�@�.H�#�� �Q�n�Q�0�4*~��5g/�E�����s�^T�5���t[=��.��Wo6]�d��OIf>�����v�����\�_�/͜�c͒����˙CNwq�e�wj�Nљ�q:7Ϗ8q���|����h��IP�hÁ���#�v��]��"�P8����zkF;����9�a��,y.����bg�lƂm[��x(rR4��r��n��H�ˌ���YT��T�n�"��$~�GJ ϕo~��*�+(vc��RI񮷫�H��D@M�@�R	� �L*���ǈǝ�%��ԅ�/}R�8/���e��cd�#�S]��uH���E+N�Cf�0h����HTlE� FJ�ɼ�9�����*&V�� 2��,2}�a�):�Ռ�	��֫X42�5kΒ����#�֩<��M�d6��(�D���x�6E�nkFc����F�c�Et=s��:������޻_�CŅ��C#�w�R'��\YB���LZQ>���;Î���gq΢?�dPT�B��$/����5�v���/��C�ϰ�+d��(�B� De�T���II a����\�1�b�s���y���N�e�|�J P�M�|�a�9/ǣ(;JC��U����,�Y�97I�ET�+�"��+�����ʫ{�C������W��݂�^�MM�F��,��O?�\6��	�D�����tV�mJ�&>4;x�|���\�mv����~G�l0ފ�Y�)|���7_>���;ѨNK�uA�h�m�ib�4#�������E#HgR0��ȑgD�T�k��0l�:u-���t��t�j5E���=���Q����� ���4(v-���f����Ze'�謆}��8^ϡ�uá��swD���#�i�
|�nJ0ߖ�F>:@B��[����2���k����>��%��B|3�����Z)�f��������4T�i��B�Q� ���徣�>k k����;�E��֯��P?��@�~3йy~����kg�<<:*BkZ:��|婭�s|��-�2,0�v�u�EPH*E������;J�X�Z��Vј� g�ʶ���j�/��̯���[1?3��{N����H�-�}$�+Z	r�e���"��7MZ��hhWk$J+֠�o ��U).4=D�+�J��Q�

�"7��S#V�&�H��	�������<VvGX���RW��h
�Mv6�^���B�DƲq��kѨT%�����ܼX��<~�P�B�{�-�l�Y)�]U,K���H4'�� D::1RQ�r��mbxx1���wadY	_�£xv����<����Z�c�E0+#�[gG�S������a�.3�&�e}L�GКK���?|?~�=�$������Ug�����/l�S277+0���c�O�LR�K���
�������Jâ2)��Vҥ @H�2Xxs�,lY����@�V���/ҡ�^�F%�&ҕ�He�������^
�Baal�B7;+���ݻw��8��+�B��7� ��E`��Fvv8�$4��t��@����h���Q��u.�s;�6u�@�cbQ�c;ळ����W��k��q�������細c�<�]^?L$gg�G���/X �VRt�.��d3Й�N�Sbe-��)&z�!��)�՟��^܍��^̜:�b!��˖��-5Lg�B�3�4�&�aD�Z������s�R����B���읩���r�ga�O �E��pDBxe�=<��,Ke�-P�����.~���l8��օ�L�-;���z����.��\��"E�l#�u�������Z�"�(����M/��g_�#�?;߃&u7t�k��.B}�3d��TI����� �!��%#�fع}�t85�v������/���q�9��������tn�����Ow����
�� ��+c�x����?р��vBxN!�;;��-U��!��`��m��BHMݛ�FCֱ�?�t��>�M��DRx������ؔJǄ�.iR�J��\�0R�*�#R�b��0.�cx��%��"�/W����B���|ī�����X�!��E���'<M� ƮG�M�O|OҸ���JL=�H�e�/���ܺ�#�����n��/��];��˯Įݻѿx�����.ԭ���|�R��x%�yr��N����� Y@ٶ8|�����kg�5��y�a�&g����i�j�\�n��s��*��P�<Ձ2� ��/���^�W���ׇ��H�#�2�v��Y�w?x?V�0���9�>���Sц����lF
h���  P�*!�] e?j-Й���K��_i=�X+I��h'����W_-���Y�3׃��{Ņ��Ó��A��!u!t�"����D[�9N���xp|���W^)`� �~.ф����$�v~�A�<�	P`ׇ�w�K�٠�>щD�=,�����K�c!�It0�#n���@/���*�{�*�^�Z�³��F�y8zlϽ��:�*M�Z��R1�' ��	�)��; �3�C��F@m(���i"Ŏ� (��"��?��o��U&s�pj���JX�tD���Ѡd�0iZ1�By������ � ��G���E.��\.#� �7�HIe��P4L��R�(�"����%ءI)�V.�T��R3ӧ�t����?���̇9�����A� bWz/q�5�24���a��Ra��|�,��_���p��˴Ƕ�x�.,h��?����klٵ����)�\k��D����2���/R���_6���atw�a��m�\v��[�����0�ӡ;U�yuG��������< �Z>{����g`��c��� �zۅ��8:�
֮�sh�q�r)Bg�5�&@��R�&1ّ8ei�� ;��B�%Bk�;�ų�=}�#\qŕ&�m�wnz!+u4��*���y?W=eś���_▆�%K�7�D�ij�*Z�^�e(u*#D�é��W��$񀥎W��[u�]j��=gE����E���+Xl�&$ =l%/A,�#I'I�u�a�ϡ96�޳V�����ga��f�e�=�Y�D� E��<D��/ ��fL�Ų�||&v���e��-9/��.)��FF�$P�Ů����'�O4����zv�\e��s��aܲ^�� �",��_K��y�{�P����­7^��C�l=z0����YI�8qJ���bo���I#P��hb�pn
�<
�\Ve�X���,���ώW�	DX���fF�&�`1����Bp�� �K�Z� &��{�t>�ߑ��$�;��.�����<g!o�����66n�(����h]�iZE�vU�8&����1p�b5��ٙ���7�� �`����'���?�ܽN�����X<�]�d^����a\��x�*F����\���2���g+8xp������]���!��V�6B�f�?�г������f�3���m�I[�S��"�, ��A��}(�N�Tȋ����C�R�R(�����|^����L���)�P�@�s
E4�8~9mW27z�$�6���r8�5"�ҶQB�@�*�v���y�k�0d��6�B;��ф��U>�x1�=��94��,�������ހ��}��R�n[���|�c���l��K�(W�2��i����s[h�
�f�9,]�y���B��p�� �������Z����:5ԏ�[���_���<�(g�s�?����|	5�������;���<|���m�A�?�e�=�ʻ��q`��}�xĂ��!���J9W�$�B�]H��=�M�uN��o������̌ʸ����*�}`�N����wj\�S���4�z�l7���,�f[�PC"1͢܎;�|(�yb�\��G�K��KL�sZ�1D��GE�g" ��HH�6�v
C�0~�(��y)J�"�Ǐ㚻߄ˮ��|�8~�4�i�j�Th^�W���x��q�V&�M�*1Y����H�S�+��Ƙ�!�l��ЏD�b0�P��B8������P ��㉠����e�?���P�vχ���a� �B�ğ���?��V���ĉc¹g���P�����ziGvJ��U�c
)r�}� $q�Jr^���tءx饗�ʖ�e�;7�6m�P@v!�@�x@�s9�Y�瘎��x    IDAT�A�<�����o�4����rgv@$>���N�"=s�z�ܹs�V�������e�]&��I�)b"H޻W�� 檫���yLBym�p���8�������gN�)YI����o�����ƺs���K.@W�	N��_����cc�����p�s�"�$#`���]�H��@�fgD�1в�5���gi��5ɝ�z�Yŧ>�[X�����}bzP�f�' �$-*0@��G��[���
�i+ �n�%|���5�xmX�\O�AǮ��!��Uq|tL�z{��r�r�;"�!͏)�-�s|�Ja*��k֠ԕ�L����
��_�A/�Z����iW=��B`�tb�G�S�D�L �+�>-	|����'?�an(9%�P(���;|�K�7�X4�ӳU8tΣ�K!43>�ݐ�D�K��Q�v�ݻ�]t�SX=<�_�>��C�U��W_ҩ�~�o�Λ:3��3йy:WEgΘ怜��F.�A�^G��0��D�ct�����1���	@H�"�s�QAb_�T��U�!�R/�*�W�M�b�X��%+�RB�r)xI���1+
��Ֆ��\Qe��|q� �GFF��Qm*ZS��|PL�a�MLUJ�� =s'�@ɔ	���؞7�_$�O,Q���چ!�Bʇ��I�0L��:T��8��e)�A[ִ�����IlM���`�\V���t:{D��`$����d��@L^��ԓ��Jh�
N�b3�A���W��0�ʤ����<�*�/�$w�4;�/p�j�n�&!r,�Hw�u����5QH�8w�r|􃿏�8_۱swT�g*x 1Ӝ'&&�XgqM�0�X33�BK�J=W�9�D�!��8�^��%���?)R^x���w�����3B ��O�y��(������W�P�b�T'���&D�ߢHR��-y衇��'� `a"рpLb�w�~��� �]��V(gV�/�°{C7�m۶I��G];DK�=���O�1ԇ��/���=/;AS���$b{���z�!���D�l�[�k`r�8�9-W����}�9>��9¶��ޭD�v��.;q@��A��G�_>�%f�������C{�(*s�(�sB�PP�Oj�6[Ʃ�	g�^	;��NAu�V�7v����An���L���E�p��<����5�ʕg!�Ұo߫0}}=�I�؉�8zlL��UkVc���h���G��_P��1���~E�*��Bi�����h1�`'&R#l[�>���෪����V��A#�8?d߁�����^~� "�fJh�C�n$�\�!�h�|���|����I�ߺe�tL�(�%�V���C�Z��ۮYߩ�:Dg~���<?��u>��9���E�ӰM�L�63��,|ቭزwN��+���W���E�-��@#qD���|$��ؚV��#I�&����]4�7|M@S"��VTB�H���K�!�ZԠHZ8I?�d�V�S(��H]�T!J^9�a� N;X�XH.��X���d�X_�?}���t��[���L�#�֙�N ;#Ԅ��%���H��0]{�9�ZW���^�=��۷�:;3�Q�8A�
��F �%s�� �r���  "X��N� ��J�@�#�jG��7�����9ồ�&I�72҆�saV/����AMhL�O��b�MX��Fm
��s��Z�yqBc�+�<L�G�� ���d�X�JA\���j
Ha�. �b�X�X����s#��#W��8Lp� �_���{^������կ
5�� 87����m��4��9%mJ��^X�4$�Y��z�t0x\�@���� �|�K_Z�)��p��q�ҩ8�n�t0�{|�k_�sJ F�D ¹����C�?��%]%��c�:ۂ�2�l�m�86z�K��-��۠����T��3D�L�&�5j�b�
���`�*��3�ѝ��.u �G
��̳���p���|����Ѐ3{��S���Eoo� n�Q�bi����Q��fd�_|�X�q��o9���N�g��%�F�Z�̍Hg�R�SOn�o0r޹�"�����a`�]�y�59:��r](�}�H��hji��w���0��e�9<n�Wa�3Azɼ��4���O�� �W�l����,�O�µk��~���rT���0ҫ�Gі=���_|7o�������!B�:�L���ٖhbl=�٫W�����-;�&Ҧ���_����v�M��n���N��Y
t��'0���'0ɝ]�vf`���hz�,�Z��Lc���KOmǖ���"n��_ج�E|�+R�,�(b7,�W�^p�*�]��ߤ��+�'Ɯ�d�������+Ѯ�dj)�I�`���B��rOV� �.��r �:�C�.��4bN�!W��ϛ����n�	gt���(�LP#+�"�P�,��^#V���F��<�z������qۨ�j*g"�d�v:&	��g ����F��c����p� D�J8�1{"^�����(�A�ՔN�s��r�h�,V ��\�|I8�x�2G%@�$ˁ�`�#��](�	@���  a����s���@��&,�  �0�������$���SP�`A��fŎiPk���+�pA�-��Ɛ����A��B�E.�sG-;,�W�p<	��`��& ����H���~� 5�U��vQx�t�b���G�����rlMI���sN8�&��m߾]�@���������\��׿�u�G���R8�-�)sWȔp��2Y�XZ0-CRƋ�.Y�P)�J?Ż��2HTCdf�$ �O"�	� �����;tQc��!�M�!����_��3sSc^�����`�ť��Ç����q1$����D�ǐ�`в��:mW�-��"�5v4ӆ���)<�i3�/ǥ�7Ű��&
�����F��� ��H�(���}
����L4��^�c��K�h�@���5$`>v�^qL����gĞ���|��H��F���&����sVc��8�L=�=x���G��O�YEx�	3�@����$�P�)y���c���r�ض�˜&��w6�q��P�H�u�r��N���z��gl:7���	��;/�r ���a1a���f���
���v�>6#�g!�d0��Q��*��Ż�@�Q�W��8$�^���
C~�F��`�!W����Ӗ�^�K�6m2z��]�^�*���\5��S�>B�"Kz:#�}F*+�%Yh5ca2)Ng�@~���]a�-Rx� ����.XT�3D�,V8g�6�)%`w0�P�������7<	Md烅�� Q !>>�J*;^�nY�9Wǩ~F�G ���hV�^��G�c� 9~��2�z����Z���n�v|m�+v�%8(�X���S=H���l��r�&��0'�  �؆��y�al�,�mqh�	���dz��yH��H�n�^�J�I�)X�=l�Ԋp��{�V�U\�R����y�f)��5 x � ��W�"ݛ$���)畟��I%#@�X�;v2���o��N�ƫ����z�m�<��cB��g	��ѡf��љ���DJ�OZ���u#��֭[p$	�w�}���
�v���u�99���VY������\Ot�s�U{�u��6|�1�3�v`��%a��a�HJ��-ᛱ�����:��>��_q>���n��/���144���E"Zg����ȖB�\���Bs\�b��
!����虶2��BP�Kw�Nu�|Z�4�>�cG��� ��]]%�29�
|����j����l��"��,=ɡ��xf�	|�s�D�A9��1,.�| ��#��ӱ�5� IK% �4Kume!!@&���q6��>7��g���������嚵�Yt��;����'7�н�f�':��.U �M�3&,3���u�`��W�nq�ul8�,����Aޯ ���ƫ:5�O�+�����tn�������?/�>��L���c@���O���蜋&�$��1�' $��P�¤�A��oD��I^^��/V���%�v�q���IHq[�2\�NF��G����oW �BV�&J"4.���'�ʂ��TV@H���_Z��Ä:tz>E�p�+�8$:�3;"gy��@��i��i-��3HX�m->6��� ���w$P�c!"��t�BT��Q��L��'�&��ޘ���`TP�jA�'�/�CH��|q�n>�	*E����@x4��Ċ�A���U��ĥ�Ǔ���"��2F&�K$���וG:����Z�-:~�E�2/`fh�R)�}ߓ♿��KP\�d��[����HN�i�� �@VK�~�� �����_/����������
� �������>�S�B(��,	-,I&O 	}���Ȏ��\s�����6(�f'�ӟ�� �~��
�Y �	x8�$L�ۢ��b��:�c山��mq�<3�hI���s�y[@�ݡX�F$l)�w���ԥ��W�ym��R�0XhJ���.L�q�@Z �2�Ī��� .nX@&p�e��'�+��!�IL����^��8"J�xH�^k�k8�0����y"6�|��E�n�Ƞ^�K��o` �C�� U�s����t��8�h�̔ �W�ܐB�^�!����c��sxf�	|�O�n.]���%����:  D:?�CuDb=W�>�"�i��zemn�!�[�}�S`����I�3LL���ؼm'�B�]}h:!����UX9K�ל��l�v� bi.Y����
 �*���:5ԏ�k���_���<� '�s�?�l�w$��֔����C:��ÉZ�r+D���o�=zd)�|F&}"�&��<��;�c4���|z��P,����Wb>��ݔ�UB��pHx�I����qe�Ʈ:0Bbp�M?�<|�� E�W��l�3g( I�-���f���[ Du5bmE\�'�nUpQgaHq���	@�⟿�P�Ŝ�.�NAB@K�@ ��_!�鲨W�6ν��b����#��: ��w���`D��D��U������H����V92؏�[�*�?��y#B�a�	� c/Ӧ���ݘ����*�F��@|�r(t����VN=#�Q*���H���J4��E"��"<t<�Ħ6��
�mЮ��
�6l�[� 97�-�8����}��'��p�/vQj�/vX�����5�E�WBc�ܓ�E��w�����#��F�`�@� �����Xt�z��e? <V��Ա$[�4�/|��?�44vu�8<v��c��P� ��ty�-�N[�&�����G���@��T!�h���w��|��lxz�\��"��t�(,��!M�"H	�����B����U����݇�v3�1�x�Jݢ_`��>+�	P�0�R@x���2�,�Vn;��t�.m�ax�0���k
���{qZ�g��V�?r�t=tu����Z��PiTQnk�����?���n�-�B��Lv6�v%yL�Hb�M�9;Ê�E�&Ա�^۶�pێʗi7�6��e|����j4�[�:4<��=�8�Γ=q
u�h�� =�\�[C6��`_/��}���em�_x~����q�5f�[���P?�Wk�]�����<���3g����ǣ�rE�bO����Ƿ���7�>� =%:�Y���$\
e�;U@K:���
/��iwۿJ�8���a1`P�'�h:����#��H	#��9I���)],l�{"�Ԟ���ą���f�z�I�BK� �U��y&���@="��P���x%����KE�>C�	�Y�H���0��9U��o��*� �ꀸmeW��$?��Q���X�/�d�<J���U4)��<�2�BjnCV�ٍ�"���P���+��3"�;����y�eɍ���P �V�&p��㎛�EJ�ᴪ��2���bpjz�������G�>W�G�������D[���v����GJ��U�B�+��|H�Kq6Ǣ���{�G �����XIH��H!OP�;,��sn���~6q���8&���*P���� 8 �`ǃz��G�
� p"���@�T2ҡ�a��}p{Q�����?��8V;��N���`�W:č)��V��/dҲ����˱n�9�TgP�����1�N�jK:#�A��©�x^��U��g�t@�墤�D�X���RQ���8�ٚr��cx�5����{��^��1��f1�t1z�d�C:����a��,f'�P�k6�h�t��#�ɓ�س�U���U���ru�K�t�b� _��m�����oLS��H�t�]@�tAB}?�s�E!��o<{��ⓘӗ��{��I�1�0e(! $�jq�B����]\����I�?^ˁF`���sDY�f����_��_r�gj��9wQJ������_�E�'�D�	a�᎖���\�|	�v�3�b��MW^���Fm\D�w�pe���T��g�s����������T ���)�#�3<�ܫز��W�l���n�
�NQa!�n�-A�,�W=	$��A���0+�����`�0y�|��۰(
�p����I�C�����5^�g���:@t�⺬ʼ����L�M@/dĆR\��ىւ�W_���G��wB�J
�3; ɻ����d�*/0�̰� �hj��n��
'����i��|OѨR�՞�����`v�u��{��s2�Lz!$��PC ��`YEW]�׊����V]몫���u�� "U �!=���dz�����~�=aP��?T��<�L������s�����[�$t~�}c?��RHB�6�$s�f	��"M��t*���I�K�B ���v�# ���7Q^H�db>����w������'�뮻-͍�����"�2]��"�E;s��U4G�D�v��' a'� ��;�P����tn�]vHq"��@�E`���k	TB8����	������S¹�Uԭ�\��<�'�!Ō�!� ��6��e�%�6A������#��8|._�"������o,�	V8G �n���~�k��_�9i�ge?����K/�s���w��>���>�K5t�ۏ������\�9)ض
��xu "�=u
V,�	; u�t�슀mS$ݙ8�Ϙ�/}���F���8���ڨ]h�v,E�oA
�(MTpx�!T�aJ6�C���x&�ay����vU�,̤fv�#�K!���s,I��}f��b|��},f�b�f�h��`�������7?�j��^
��M4�~�@���YMH�)	3;x��!��Z���f�*�e1�ӕ"NX<��M8����s�����ǟ݅�?�qz�T��@@��k�dRY�ڹ5�E���ʳO�%矆`� RJ篝 ����Q�9f`
��9fyj/�x�������~�D�,�{6b{�lߔ�_7L��]��ep ?�(`�>���k�0��v���~�Rt,*
�1�B2����z �5��T����2)�r�?�#ּ5�Umy��|Մ��ER"<�#ї�̆���#�+1z��WH�R��[���.}^�?�#"Pu��H�^G�9�ܱ"0�hF"SIk�bM>X�L�|IGe���K�iA�CP(�41������ԳA&[�3����"~+��{]{B���Hv�|���jgҦ����P�:H�ڼ�2������
梍h*���Sx�����ɟ��g��۱z�j	{caNw(��	X\xDZ�d�U4�, Y��`'�-bcf���E �?G��,�#�>���ц���Q����n��o���$���&`&��nC""+>?��N-�9ݳ{Ap�G�"�$	׉�1�/������9��x�~E��@#+�9����7a������w��7c�n��ر{�ش	{F��Z`�i؎
��C�y�f��-���3POD���k\�g���6r ��9@[O    IDAT�ׯ{7����=8�{�3��7�M��̸>=���q�U�B�Fm���D�x
q�]W���=��ؖG�H)����G�!���8z{B!�.�w�P4_tg���\c�8@�L �J!�k@��q�}��[ףh�B	"��� ���>�����c�$�,���@�1�\b� �J3(�C��RU�mH!����q���_������ N�?S���{v��C*��S�c �3f�1ۂ��w�{n��pѹ��S��Q�A�n�e�M%�Oz���qj����v�֦�<5/�ظmw@�
_��,5& �?�8��(��q�rlv4�N�+�>�
���X��J7�\��!�9�+�k>f�lA\��}ɤ.�ةdLl]-Za�ᇪ��8����X�Q,�0<4����r4��oM5��iJ���i$m��7���0�O�n�X��F��*9���֥su����@~��otY�TD $	�]��I�[/4�:E*;O�uIw�	)2^څ֩2�dr�;��10����c��߽�'*�*|҈���[B�Z8��yp��:�1����<S}��g>�x��=�̵�'�\�/�c�q�bqL B0@(v3XXG �]�� ����D4�(�"�L��Q�����
�΄���|�菺'Q�xT�s�|.�"�c��Q�&���B}MhqM`uh��An��3vi����E{^ҸxL�6"��i9:8�Ȯ�se}D�+�L��S�M�^_C���[p0��.��ކ'T.��[�㱧���!vX��� Q��s ��+�qE���B!+*��!�g\.P�H�ʃݸ���ʧ߅x���#���������t�r�������v��ij�\�<N��
��T)�s�l��7���Gz\�L��ÒyR)U0c�L� �X�{�(Q�<��i$�)h�=ab�V����A���A��oȱ�S$� �؍��:eɂ���^����c��<�8����8aI'����ߋ]���_�:n���&8j�+U]s�"�Њg7o��T�!�sN]���:��>��T�y��?x���?��?5���y�dS;���<�쎠Ƅs% �&���}n9�Ƿ��8<r�K�0��)a"�$�ʫ��R �(�ap�2� �P9�͘;������At�؂x\A,�"�j0i�[���9�,x��OyCc��/��apt#�UTj
U�Pr�I��,ۇ�C� �`�j�̷p�LZ,��R�,�=NR�D���Φ���P��|��o�ґ��w���c"�߲�ZSH1�:!0y����#��?׭�s����]ǨZ�@���_uo����Q��e�a��D�`
tM]�Y<��w��$���	&,��|d3Y�=y�TSEc&�K/� ���efv��,Z8�y�������$�"���u��>]V���D����+�ED�'ҁD]���e+& � �N�+ �Ŭ�\�!�+*��w������׈�,ӆ! ��pG������h<ѹ�4!(!�!0�W
�mvzh����p|}�-�Ec�:"|.�ñG��E�u}��(Ä���J�MX�|���!�mUVq�lz
��a��xz�����H@zR�ċ9|/	; ��f�2 ��×� �N�֠yL�OGq�W�j5��×�,�3~�}G|�E�Ď�nơ�1h��D��j�h���Z5Ԟ1%�4O:������_xu=��'��ۏ=;�`h`��fqK%Sґt�j���j��(�C7ݵ߻}=��y��y��V�[�G#�]\���|¼��KtY��=1�����
׆�Jî��H�`��̖\��k0�kFG��ւ#�����Oo��/d�Ì3�K7c��h�6I��ůX�Ջg � ��(X/���1�hf`
��hN��@^3�i�^��c����z
6�޸��@�cR�����V�C�1�:�ff���JWD#%�)"�0�)�UKg"��TFq�¹hJ%�x��¥{"���Cc6')�aA	TjU���G7>��z�g�!CCS=��c`p����e.�\ua����D�

�م��-����H$��c&_���#��d Y�YOE�Z���D��u#�#�|��yM����'�N�"�]��B�^[�nD���+�Ѿ&oz28���c���#ږt|xbX;Je]�.��.�[�qƩk0�ߋ�{�ѷs7j��R,��\u�"&�����`�F|�ס1�D_�A45�0:2�.��$յ
{�wI�=c�,�CuwwK1�)"�t���s[,��u#��xN��k�4C��\$H��i�N��c'�E}�E�{T�m���Ȳ���_|�J�KD�" �":U4ד�	���lu�/�?�D�帢}F]��㏜������u��D���]����Iܻ�4���������y����
���w�=�8:4�2)�̘�t�˼v����)4� ŉ�qɺ�d��8XIאᗎ�gj�������g��W]el7�B/F�oʡ���I�5f�����Џx��S .|�vS�4�Z�"��܎7@m
�¶$̔X]�e�?k��E��2C;q� *S�}媃X<�@W�7a�{�=�o{��<ر��4	�0�Hn�z�Q�E�@�s�R�ޘ���\�c-�^��&��$���*��-�i'��?^���̢�O<كO_���l(F\��t�G6��3��J��E�'���ii��hM�8�)
֋�s{j/�� /��65�?��>��O�"��x�AAI��va��}��,/�S���t����5~͂��H�L8V~��T�EGK���hi�lN3�t�0��3Z�Pj�<���AT�E)J	dU�i�*͠/Z�Θ=J"�r�{t��[��|-�ln<%�����++��+�j�A�!�A<�D,<Xq�;#��������`T���{�U�0?�u=�q��ѝ"M� �tԻ�����Z��������'wW�"rrGd����uf�5�=�I��2ֺ�F(-t�aW �"a L@��:5J!�.�UEcc眽��Ȏ]�eon�R����WU&�ڡtL�駜�O|����0:�C�~DCQ.�����7
�j��nL&0w�I�S��.C4�HR�YǨY��B}�I�ᴐ��%-[�!�#c  `�t�D"U���V����F4�Q�!�,E Q4Mu�N�}>���_;]��?GnTQw$Ҵ�;_˱s��߹}R�"�=)ZQ���GD/�lz9>�/�;">�&w��<����p���&�������+�	�����R���bOK�B����jH��'j��i����&���7R�|&�����<��"xC;�r?��F��҈Ɩ�8.h����Lz]ԻSqY��!��fH�"(�I��L���@: �Sb�����0����X̔@O6=�J���bœCO �I(92V�?����'PḾ�7�,�{��6�2��K�GX�H@c�C��� �t�餧H$�([�Y��H#5��U�kUP��ɧ�ƺ3Oǡ�=xz�nt�끙�I8�M����D�}v;<_�¹]8��1F��(b^�}�T�'�,���_�L�<��x���880���KX?�5Î��7ĝ?�@K�j���5���
�|`
�G\g���2
�-`��K���Дp0-�늋�2]{�k�f�E��'��-�x��qY%��+�ɤ�X"��;�>s��
�į�=GƐL�!�s(�T�U1Zr14Q�8iYj~�₫�|Z3lD#E�U�%�@,��J�Z���*#]a��+�1�ƤT�0[]��N��=���HP��<���s%f
����wpl��rZ'�����~G���6��F�s�x�ԝ��)S5]\�X�1�Y�V�T�SC��0z�T�&]���-m�Y��,��S�Ij8��SМO�V) ^��J�?8�]�v����b;4�/��3w��_p�X�DŸ�3:��y�昦H׶�[�k��c�6�L<�z^J�a����,���t=5<�΍ܢ��`�B5�C��r;,�# 	��^���?G]�-.��5Y\�1q<|DY$�8>z��>���[�1�+�dZԻB$�wE]�BՓ�y�|�t'��C��)(��b|l��?P0ɷ�8B��3 TE��91`џB��W� D,wDH
V6ء_��%��"�H(
J��p��_�����p�C��016���&4651,�W�����U�� �p<�4ǠK;��_?�	)��TL(\�JE��MZ(:7�#�x{��1s�=C�&�q�̔dլW�[�MwoB%щ��G�6�$ 	/��=�`Ah� bu�������!�[��<�m�q��'h�4�2�8��r��\cfu�@s�O>�����ů<'/�B֛@"(��u'O�P��7��L����g겘��I3���P�?<"�f����AK��>��{���L�\�E�Xt��$��s|$�2:�\x�rL�x�l6q��hJjص�i�ٱ-�s�l��	S�Y�䳍���ZUR�+���V��豸h<�,^��֮Eo� |`#��Ө�1��30X�1V��;Z��Hv`�*��S�!|z&p���cI�,��8�αQ�&B�/�u�B��p$�;E\��HqѺ~[�N �!�I�B'��f$��w���~�o�Ѿ&�ywB�z�$���1IZ'�d��br~�"Z:
j㢬'4��;����S�zժ�f����I�U��U`�t*�Q -MM��	YY���𤲑RAלyb'+S����N���m*\�W�#
��ۋhk"4�������7�ՠ]-�f�HH����'~���W�3R*K�t�_���N��HG�dq�+����=�G��|A�B��1Q��c�}u>"*�A�`�v��o���`�A�ϵh\� �T#E��R- �M���5�B"�|
�lJ��tB4��Z�WK�� �5��1 "�(�+R�<f�I�4�����q��/C��6Ľ����ۑm�C5u؁%ZgČܚ�D<��2|���8�f�޽�^4}z;<�G"�X(UK�'G�x��#���v�i��Ù��j��P����2��Y����'w?�Z2Ԁ���N���\D:t�{rr�
Ay�d.�
�]�E�|�!���!xt��q��	S�iI���y�G�r`�Ң�h.��H7�ǒ�_��dF ^���q���HY#ș>�9}�T5UAL���r�n����M��sv:*I�,���<=�������xz�Q�F�8���ʼ�UH�-�^�?���NX؂ei���'����R�~�밋hmjD&���p�Wĳ�L�APta+�Ò)֦��(rv�u�XE�qpօ�D�¥��ǝ�ݍ[� ,$`f[Q�u�Tp��8�5������n��$`�b4�E���P��H"Й���O͈����c��T���b�!,>Ę���:�GrŞ�X#�[E�,@�숗���B]O����9�?���:xRX�s�F�kX��QW���%��=��	MB�Nz;d�ŁJ�������dL�I
��L��DW4�P�$�e^�L�x���f�.���;O,���n�'`j�P�XX�9!P ��# " liiłE�z�J��p�g��[�l�a��6��E��vGF�p����B:S��ϣ!ժ��L�f:zOO���a���}ttX�
;5d��`��3���ZM��C�A@��7	����q^��	V"�����n����R	�b	)D{{�仄�9��c$����YptɊ�7�yi�Z[[%� ��o`#�����+Y�n"���w�@���Mj#�,f���>�JM�Q4�+a��*-_C�M@H��98��M���CL���^���^��\~�G�Ȣ��`ftLG��	:�φ���TI&��H%�s��BE�?�j(�?�o?�ϛ����n,��[�2Џ�S�	h���$����Q�W�{]�%���	
*��1K�~�7ݽ��l��&����c�J��Ps��&X����σ(�B�\������bB�����5C ����>8���<�]�H$����I�|U�?3 SA�0�k6�i�&z�c፯}�X�^i��Y��0UC�u�SG�g������0�S�x���ֽ����I��$�������j?Xu�v�$as��.�	U$�A�b�qX���P7>v�����;�]�6�@��L���j?�E?~�ſN�U�*�["fJ1Ă'3�!K!qi��6_g�p��5Py|��n��Zf�h��7l�w���Hv�ENR,2�j�B
WԍQ��HH>H`�0���:�����-W��H�*<��r����6���r�&+��d�cK4���|V�=�FB7� G�0��[F&ۀRH44�jSG���b��"�X�!�D*-Sρ����Ȥ�as�=:#�A*�ge��r�D��bj2�v�;$�1F<��<˪�Hġ(T-@�\�WCC�q����.䖋����0�����mo��U,_���`3�CGPcv�)�=Bc��$�N�
�6��\LFalT�(�}I�c�Yߎ��IWa�%hjm�s2Q*�y!`!O�Nd�K0<�(8s�t),ҹ�?00 ���t2t�J���:Ӧ�aZ�`��R�wvv�u�{�n<��3�y��aƌ�ؾ}�t*��Np��߲l�Aŭ��*7Xx*� �U�N:��E��AI%�s,V�^݉�,B�w��͛� �C��;:�biB�'
cR�R��}rbᛡv����±s~��M�-���s��rU
U�Vܢ�p���W�
���j����4�B]55%5G��|�^�`���:|�"}]lrA��<� ���4ރB�8��zk�Ƃ6ۅ#8k�4|�����>T�c�蜎t*'`��$�U�EJ��:������C� �m��1.Z� m�Mhi��H f�m<� +�{8
&����]s��Bp��AҜ�)u�J���8
�
��<�[h����&p���o�����pu:�)P����1Xt���C����2)m!x�M9��J:n¢�<C�P@��J�A:�ECC��G0�s4X��Z��Rs�g���^�6��-�3yxiH���M'1��E�Qvn�SՐ�\pΩ�`�*$�Қ�3V-���^:�S#}������";!S������G���~hj +��Î�a�������+H aA�r������8ii�^��)Kg6�I)b���q����	�u��"a$��p�X.y�����Q���C>>ݰX<6���j)@���
�$��`�38��q�o������(�-s�n�������?R�Ex_	�߂��`�<&7t�JĠ$Lht��Ǡ'ҰA�&t�T�Dq�(�	��f��Dg˅��
��z�'�
�]��M�\i��Exv�_�z����pt��x�E8���p
�gt��s�5�3f�Jx<��61<.�%�%��P��?��
��ϛ��W7`4�$P�]�L:��X)t,0�daw�(DC2��u9Gvo��I �M���L.�H�X���D�q�6�c	��\��R��`Q�ll_�� i��h�F��*"f�b�l��+�1U�]�(���h�';\��8Ē�c�vb���"� �]
�
m�Ҕ�.],��#G�`w!�,ʣ\�һ�����f:��m�,[�L�y�H�$�Xp��ǡC�(-^�X �vP��>�|�t�M�m�]Ǘn���+�w���l��bG�@)��`��i�;w��\�R����0iVԶ��/R�֯T
�Y�2���~X�>�q���r�;�����N��:-0
)����MԵd��� J�T��
�hH��)��{�Je�k�܀�,�y�PIk�ފ�6Ä�L�/�(��4�f-��D Ⱥ���Ͻ	gc{0:ދι��oh�qr�D1,��*�����?����0bi���*�t�Fk[#��$Iz܇��p�mC�`bb����aT&��f��� �`K-�n�H}    IDAT��"n�y,�sa�M��;6⻷='7U�+.�T��M��U���p1��˶�TtT+e�vY�u��X*	�4P*�L�QG��x�[ނ����%tv�@��ޥ�uOoڎ�����ݍ�=�H4������
�jF>�ZA&�����`h&v��͜v�� �y^}�Ы�h0|�ur��2�������g`�����l��3�}�/8�*�T��@w_�nڏ�6쀣6������U/�P�Yť�-�y�,�������wߊ��}������&!��T
c�t@��/��D"Y��uE�h�좫jղ$f':Ҵ�tjH�⒔�Э�b+N:�V���'6���SL�h��c�z-��18\�3���.�� ��|�ܙ�g��e���������Yhoi��/~�͜���1<��f<��S��,�;">��b]��:��&4x�Jx�ړ��/]�����ӝ8�?5��"�@	g���/}
�2a��
62&eW-h]L��������^+��~��O=��G�Bˤ`seYe[E���H6�3;$ż�ՔN��H�)`NG+N^���Covu�ǯ����p���㧶��/��x�C�t�t��єǞ�φ�$�f���k[0c
�Fy��́S+`t�(���Jq�1s6?����A�cY҅�;����g��B�}L\-t�$� T̝�%��=Ga�SOa���ct'��ȥ�E:s>�n�(�U�V	8	5'�>�Y,��<�C�6
��Z�t)-Z����g2��PԪ�����Rȳ����$�!͊�>�!�Ia����ܱc�ثV��c' 	�#!E�
������GY/��5k��2��z�)q�#nڴ���Ç�(���Uc�"�&���r@"�=��t�|qc�(��"n���T�lԤuR��x=�g�Gx���Au ��=�}0��]% a����U��fA_��}h�ڇ����3������Hwb��
��@`�nt� zj�*����&�3bW�H�
eÁ7��E��LT1pdC�r�4�F1\��aBCծ
���X�()|��G���CiZ�b����et�8�8�^l�&CU-!�N"Pjx�k_��<���:K�R�%����}8��s��^�Y��p�MU\��������.64V��[�⧷߉g��G%0�$3�B�IIw9�01��]4<;�og��o�u'��Nd �=e���+���O;S7ϟv~�����݇���@,ׅg$p`����܃�7�[ b Eo�F5$Kg�p��p�b�jJ���Mx��;%�}F��w�G僐��8�A�N����ihm��|�EVv��͠���>�8���{�V�i��Ր�)H�u$ɷV}�r`~��D��;sV��{�?��0a�N�[��H�%ãv]��o�Z*j>L�|�F�/�ԙ�f@cAR��y矁�?�.�# ����?�	�r-�<�Vb�}RMu��>�H�1T�X0o}�%X�f6<���_��G7�lh��g7�³���7�����	���\sJ�j�
]� H�#Q:�F��ش�������G2�62��:�F�R���\���A,�h��>q-�_�UԂ�+�(ό��>����SH7��7����8!'�|���E\�4 nҞ�B\��]�
����	�3jj0U�u
�y��7l~�	�67��2��j��/~y'6>�$���L:�/���E3�N���Ey�'�1�#��"|ΜN�m�����쇠�"lR�>X�<�����y��/_.wv�Z9fE%�@p.�Y`������htvv�G��Hb�
���-�)�*����� �;x\�fٶm��qٲ���iC�_��Z�X�p��8( ���yg���M�J�t�|�Q���t�ƍ���0�#Y�F��H���q�D+W���O?ӧ5#����g�F�P��}�{T���	m�qu(fRt �c1�<��%K�'��GK[�Fg2υ�$t���*���͎��|�]����a�����Ӑ���;��TX>����Mql��j��i_T$S&����(�n�/p�ϓ9`��`{�UQ+ax���[[D3��^�|(�F�z�P�_U�ދ_<q j�BLx	��!H<R��q��Q7��	�
拘ޖ��kVȱ������܈���Nh�F�?r�8T�����2���n�0,vұ���tWT��\�=�m{�bǾ#��?}�]pUM��L��)Y>I3-]���W+���k�;JiH �ygL�`��>⧆�"��) �":SC�����}����	H����c�ppۣ��tw?l%#�5t�aA���>�w�W���>���߇�	RHI��I�cY�`t.X��ǭ��"Ѽ�t��ѡ^ܻ�<�(&F�`��<�)Rl�˭Z><5#����FC����b��%`��poI�0,P��Y�P�@!5i�<�XL�BB�]vo��8֞�_��h`�0H����W�u#�F&�2�Ś#9z*#z�\D6���kރ�]p
c@�6�\kW����e�!�9v�b�����勚����(����]ŠT��1���V���=��?�/����ZZҧY��)�����!�^���t�׍σW-KJt2��x��j�b������v<��&�?؋L�9\�&u&�d��I⊸`9�2�Zp�GBq1����NZ�e��l�x���̓�O�8��ӱd���9�_�} 9bћĮ];du���=�j5;�n��E����<�;����{��
�YX���D�;<&vp�����a::�3�h>��v�#vm�ק�_�m�{ｰja(!����u��lٲM ���.]]�e��p��>v4N=�4#��ױY��Em
�G0R���&Ǔ���1bG)�La���H�Su;�P�%������"^�F瓟�4���-�;_���g���>��q
���t���3�q8���y�<@x3�G|ĠB�F�v��p�A�_D�����uX2#���U��5͍!}��@��<��@vՁ��(��)�!=Lc�.f��sCH��ֆ�<�M1t5���C6;y��щ	8�/�x�Dͩ�F-�vu�S�Z_��=�e}7��<T����&��N`B�O��*2�k�".��"��m�Ck{V�UH&�����7��֐�6ձQ��-��5W��}��g!�I�V\Ē	��#e,aĄާ�&*>�<3�k?�������2}&GǐkH�}�����;�v�9.{�
}�'�;i��/��=5��������M�{j�73�c��`�X�"�op�Ǒ��[�{J�I�m�&4qw�w$�/z�OS������_߉]pjE������ �X�	�[��]sk��	ݱ����Oc��8�o:��d��t�RقO�@��9�L�<�l��oߋ	;�hĘm��ѽ�<wZ^RHZ��ZX�:@HI���ſI1CM�j i����?�^~���ǰzf�r��o�v�����y��F+_F,�+��2NY����+q���g��ua�\s�u�.��4$�Bܖ�7��z��W��Osڳ����R��A3bHǒB�0�+�g�\ �i�t㉧�ذy~v�=xdóP�,jF"!�I�ր�m|��w�̓��)W�(O�s���=��򷍃~p��w�K_�6�x�p����Ey%��&�����7y�z��4�@U\x�YXs�b���|"N[�����<�hp�/���ܔ���+�{���'�|R�9je��G��Q�(��>9G�L�n411& ���嘍.���+V�sX��P7�N���vx����ȧ���
�LdL�����P}�����ku��0��sΑm<���ɘ\��xh��B����?&ǹf��"��P@:��	�#,�P�#��Ygh���J`$�m�����vyZ��B!?Ժ#�5\��΢t���Ў��.�Y�֢�1����J���1ttP�Ѿ}02>����l�o P�p�Ţ�Q����=).rb'~1'��+���+AuigW��"73�A*�`��V4暄1�8���X,$(�ԕ@�K���I-��}D�'�K�a{.j�#:�d,�O;�o������RI�焯%�*��7C΃��^S5#�������N8sa�9P[3��*%�R*��|ۓ�ƿ��'�ՙ��� ���i�;q�?��،�� �kFqx�}畸��P�GC&����Y�Cc�B�jl���SNj�q3��}[{�tc#�
|�'�����$rM�II7dДoq��]{B0�c� o��I�N^=UC�o>h�^35��������������q�ot� �L`�X��ߎ�
*.�,�8�ЕFw*hҊ8gE3���2؇7��_��V��魰��t<�D#$���31{չ/ȇցͷw���)545g�N$Q������(�x
�^~��߆m6b�f��7��g�s�(F�(P6%@�(�P_�+�F��E�
�]���F�d�4\���p��ʅc�	�i�)���w��םp�8<�1=�*�u��K/<�����J�ko�G>�y��_�ȴ�P����y3����m!�����~;�{�a9/��P*#a&���Q*���3N���^+9]���Gw���p��j��������������3�KW�����x���(��sd(�?�%�y��oN*�A�[�������I�~�.����e�ItԚ�݈�o>g1�?��
c
NY}���K06x�Lo|�eǮ��z$���p߽HO=��������{0>V@ww�t<hK�dDI�[,\YhXV������J�C���A�����8�H�'�R
�	8@XXsu>�+IqOp���s�cf���)�ԓ��]
�����E*j9�ZR��E�R r��l��� �իCi2,�	\"��㤦�sDP�+�ca�#)d|�u,�{��O&�R4��q�{�����-�/�m�W�x��q-�Ȧ8�o/�ꓮR__?vt��ha���5؁&]�:�1D�)@�i?R�  1S�y�F�pq�����ǐI*�=��DJ�$�c!�N�\)�uG�
AUժ�������b�@�#�0
Y��t"͐��ۚ[���A7��p���t����X�WH35�]�%V|�{�{�f��彔tM����E3��g�����>c���B��H�����r\p���*	b
�����񪵧�VƙKZ���\��O���r�>�ל{�|�e�5k�-��w���ހ�}�����&0m�y�޹K�U��ů8�[�:�|Xw��	�>A�f`j��3��B���M=sj^�3@
E�n溰�˸k�.l�G�1��	x���vZT�lYw��x���O���	n�AKPc)�4��ú7^��sAup߭�����hHƐN%A�#�'�e �Ɗ�����^����PF5����x!�נ�ƕ�I9�^b�RC���O
�@e��=w5���7���¶��m�Ɂ��AKf�p�Na���`U���s���iI+߾�����~ ��(�tkh͘���?�I󛔭�A*݀K.~36oَlc���9A���B�i�f�^v1�����8����-!5��%�9�sx��e"�N&㨌�ᵯ~%n�Ƈ�}� P�*��"�N�t,����x,�M��#ӗf�QV���"�O�eB��ʊ2)W�x����1/B�6B��	����2�VQ���d`G�+����A@<fHAN�6�#G�J���&Ј\�B�pE[�5~��_�����a�]�윍��Y4�`�B� ��=m��)2M)�Y���cq���zg �qX�d�����!!e�}>�d�N��GZ?����6M��P�7E��_C�s�v鮜r��o߾M�D1|OO���/���Gx��{����X|D��G}T:&4��<t���J�0K���y(Ҽ���E�j���8~%N9e��Z��H< �J�dO*��_�@o/���|�fhP̴h@�yaM�.4�C����k�b1�0̧qK�h�U��w\�e3��ڇW1�%'Z#:?��.&.i��+NV��u�hN� Ȕ�J��F�^҄Z��J�I)����W���0���e�0�]A��ϱQ���|���k˵�W����>�_>�A�BXZ���K�d�K�1�T#{�q��߂+�t1��>\�v�rˆ��/�Fl�~��#�k��t��W����{ax�8������x9r���.�e!f[8a�"����c��J���;\������3H�[P������,#�\��֝�y�����W�`��/�OƩ�M��?S7�?�S[|	���]{��RAB�X�б����Ѝ�=c(�4��/�|��%�b���%X=+�w�Y�%@�)�S�%�ޱKN�z�=��������<>�\Eu\YɬY,U��ox+����@Y����X-��=5�ZR$H8a�I�!ŅB{P'̸��Ơ4`���
��C���UG�w(�����+�,Ƿ�UWO?ۍ�y0�ׇLR���߅ٰ3q`�t5���_��7�J35��Z�1������NX�����qe�eW��
#�F@�K'��)���#ýX4o>�p��e��U�G�����.�烟�~7�wtbh` V����8��5����V������s�o�]�A
���?g�����
�t��>^������׀�D*ߎ���c��X��`G��2����,�����lR������>�sNY�lx�01&�1��5 �`)L�C��l>'��[��&�Z�<�8fa�2f�$wjqV�x����?��a��9�� ����#��]>����Y!���vHX�����p_����V��Cg��B�"=��'@ �x��e��Q{�mG ��温!``d߾=���Mv/��+��a�����a��t�ۖ-[d���C����"8"%�`��|0�� �_�S��#�S�*E9���6�榬tAx/��C{�0dT�O~�3��STl:���.�.D� ��59��Žʇ�S'�]P��!��^,h���w]���Ƙ�-"�2�R롨�k!0pŸ7�!�
�����]��Z��bBh���G0���P� �&I���	��*4�;6Ԧ(��%fHg'�% ���Q32��-���{�aeg���a)�d�J5�&'02����o/�%�����w`?��w���ף�e�k��}֮"fhh�g��� �Θ&�k�>\����O��2���'Xq�R\�7�aqg\.�����?��v�\3b�lb�њy;b�W�x�߼g��Y�ǩ���_��SC���Z���ej�S3��<�v�
J�J��H�[_Ŷ�q���nID/Y\�6�Z��c^[�:m���U����Z�>,�3t!�mdC-]X�d%�s־��[udK02��GHС=Q�R�.|�WJ��o���C����M� A|:�+��a�P�B��$@iB?#�T~����P�/&$bq�L�F�qښE���_?vl;����Ӧ)���W���p#.��b\}Օ8c�LeG�@����՚S��9�u���llC�F�(]t	f5��_� �d�W_I�7\�g6n���CI$�V-qb���9bO�:%�<n���/aAc�{\~�g�_>�(jn������z'֝��IE��;�[��aɌf�_�{k���C�f�l������ݽ=��4�*�#N�O~?�Ž��pe���V�e�+�R�	 Q$՞A�hS)�xښӢ�� �x�:�:u�O?�46<�Q
mױ$��]�����Ƕ��VCd��6��yf�<�G=;����O��_�0���9,�2�B�`#Ljw��_0�ж�H�"E�]	
>�gp!�
�L&+�,R����%�4�Pf��t3�R�Z����0L9.��V������ �1p>��!]��(�S�y�!�R�Qq�%    IDAT$O�!t��uنА�@���:	I��X�4�I�06�֦|'L_g'��`2�GC�J����P�",YPbI���>��1����<���8z�����\ToC�� �Z�hm��kvء�kV��\���B�'IY���B*�2�z����x�j��x�r�|����=��`H#��a�:3�� �����k�M5�?��m��8V</9 �B��Ѝ���!�Q�4|�����Kq��^|�߿���ށ��.T�,Iq-!�ˠR��~����a��#r�FK6^��k�'S"�O�L�M�$F��鏾�=���x���7��w<��G"�ǌP<[�1ϱS���7]��+"퍢Aspƚ5/�{������f�%2S7�K�DM��3On�& D�nASQ�l�ï���kχV��	]9\r�"\�W+_���VCC� ��F��J>�9K����k���/��6ܷ5Ђ��0�<��F\c`�:Ҹ��\�ū��}��=�0�]��Ş���������U]vA�`c�v'�ˠRT7�Z�NU��\�3���Sx�+օݍ�����E��-́���K�n�\�_wO���]��S	���p���1Q���1�kUq����՚³w���X�	��oށ�6u#�k���K�sPh�[)���9ǭ�9��~��0;���~���|�����x����ׇ�����ܤ����|�Sزu��;������o}#^w�+p��ٿs?�/7_���T=�Vƚ��a���B���e�֥�ͯ�Pj��Zq���,�ۧ���xAnv
��U�f���+�Y�`.�C�]C
`� fL��Q�.�Z��A�P�b1�bE���,\�X��М�� ��G�n��T*n�+�*|p<,�i+Mp��q�|>�d@'���g���K;U�D8�h����� �����&&�L���#������i��.)X<v�$%���(�<Er��;Q*��Dt�D�Z�΄m��w��'(�����݄�@UbplE: ����$Z�R$~,����x�� Hy�0.�d����ly�t���-9�Nh��LO�|&��8�]	dw9P5&C/�
U)��v�x­��;���Q΍U�7�aqn1[�NY|���hUE�BS	3��t��g��6<�k~�|��4l�<� �X��B5��ޘ�G��/����~\��Ŧ]���1C�U�[�Z%��@ܱ���w�]o~��Ў���{q�G>פ؟6�.4�Bc:!I������3W�R���t~r�C���&�^8׻w���kUq�.��+"�!��Xw�/�{���nj/S3𗟁���/�F�"��'7o��*HY��n�ad�z��FFVG)R6�1��|&�^юמ6���e��w�W �ڌXk;��9���I��6�RD��pp�6lz�1ɝ�`2����}��4^����7����8Z`p�6��>:
��Ũ	.FC��FzJ �NNfL�#	ӣg�i"Ťe��:�U+�a�-ߕc��3��5��9�i���ǵ����[��!�fL�8Ԡ:l�8E�jO���Z��CcAgK^Y���}j'b�V�:����^C&�;R���U��Y��֗��Y�?(|�ƛ��|������Ї��ם��	�Z�fv*���g�+�9����!��I�0�6Q,��o�p���oü�&e��=���X�ѥ���o_�ⷑ�X�Jͅ�.��Cz{��M�^
m��=�a��Xu�ȦT��A�]�NU
u�$�DY겈f1��ӆ:gϑ✅tX�r�>�#! ��>#S�Y��*��Ze�!�`�I0���	���!�p[�Dp�'��}�[��G�����_�Ϝ���>"�wHbw�a�J�7Hs��7my����Et0
�2i9�(��?�3I�/���� �.	��k=�:��&4�DE�s�D����1��y�E�du�1J��CSD�]#}ˌ�H�"�)X�n�uj��8Ww��>�e
���S�Ph^ ��]v���S�w�}X��(yDm�4O��s!B	���p���#]�}R�n�NF�;�X��s(���k�} ��1��^M�C(�ԋ�c��χx���hM���8{�%��4>�ݟc��h@�|Cl|:���v���U�R>�q��K�K����|���	�Ͱ�$�]�l�v�$�ϙ�����8o�RQ����'��_����ڤ��hH%P-����:s���NoR>v�m��o��D��v��eb*vl�����o|N[�@��Ҋ��N;�O��"�H�����f`����M�Ԇ_�3�i�ր!w v�`��u�ƽ�qxz������"�q�	3q�Nt�jx�׷��0�P镯 �$:OX�e'�=9�Or���j�a4���h/���: 	�N��0\(�o{'�?��N��\�9}�lO6��P#��W)�]@Q.�ؽz��"zm EQi�H�$�l�&K���gN�����?����~��xEw~�v3s��9g�}��)?���v�D/*A&*66�P�,DݧB�4��ФrV�q��x<�����2(��b>>���[�>��x��&�E��5;��;�{�~n#��gPs#8�؆ꨢ+���:�Z>k��Nx��=���E��U<'=��'21�9�l���Ob�ܬ�������ŋ���z(���>�Ȱ���g�����G��R�+��1hfO���y�p���
�=0:-�1K�כ]��O!�9O�������D��� �eH��Ɔ ��_+�6B�����	���0Tah�SI��?n�&�̂}���2q��B��:\���)�V�P���jJB^>���nɶ��V��
�S��*�[�$\Ա����>�b^�O���g"=��@:�u�\�(~��Z �5���rC �5������- ��nC��N	 !�!���E#������S�ʪ�k�`Թ���΀�3GCZ2�	u�Р�._c4t�����-�d��D���F�BM	Q(���G1����#�,jI�]& a���N���G�cV`�s�eK ,@ӿ{�ut��-č�8e�( ���=��h��	:�*�kBM���F���[�\�E��L/�z�4kU��ƀw@�<' �b�ja�7�z��Y R�2p�PܴNY���E����B�q�{ފ�^���n�x��p�}�G#��g'� ���NBCP/c�%�q��'���{�+сD��iﺎ�i0cUB?�����Ӟ�1�\8[����E�ҭ���"��%�5G��o#�dp��ן- $^F<���c���ڗ����>O��_�/JQ�����k�W��a֭��"�.r�l.���7a�� u��M�a���x��y�4�1���X��*­wu���u���)/�}�k�SQ&�jTq��o��0#�TX�e7���^�ݹ�����mЍ�Sv��B����U�<X(��*�\ia0m=D�V�|&�.xE	���5���瞤�����@�����o�:������K1$I�t)�gaa�6��oa�NK�>R���h/�ۣ������I�X�d_Y�&R	T�̟ߍ��~Vt������~8z�DGW7�s��p��fi[����{�����7���0��ۋj�&�"��Q�[vF{-���u�>�-z�>�m;'�6�u�"��IT"I �j�ꘅ�����²�a%��N�!W� 2yҕ��$s�JR�b)��))�wAa��Y�P���NGR�*�{(E8s5ĥ�Vۓ��Ɇ窢�jH`�^��"ߤ�E~V F(`���֖�����K ��3JcB ��PSC�W�h��<6n3S>��>�G0#E����[u�YD+��p����ޅ��q��ф�uq��>�@����̩N+K�E���q;|pE��|����#R�h��g@[�MLHϲc�n��p�0�*��i��7��;�{NP�m*���3��M�����_�ܖg�%��ƀ��#�;p( pkU4Z��W�b��A�T���}���2a�
�H�I��L?�P�L^g5�G(��@�<�M!�Ɋ��T�,�[��څ��z,��Y����K���ɉ/�˲c� !H0u�yۅx��"���~?��~�f�-�I��Ű�_A�,�av,-��v���> qK�|�'L\q���U�`rt]3f�{?�7}�{Hv͆��J^�X[6o �ؖL@�X��� ,��WM������}xi���Z�4�dz���W`��MQ�R�4kWw@ r�#kd�0�W] 3��q��l����:v�}�F�L�A���)�|������UMm���j���;�W��I�� ����|��_��}��xv���Yh����\��\]�Y�0%YiT�3���R�-'yZL��K�`x8����AQ�W�G?t%��Y��B@28��G?�E���������E���% (ᔓ��/���F�x=��:ι�2l�>��E�)��X�zRT�+��ς�]�����#f��ߺ�����\���|���O��)���hAg��~N�����w]��"�$�
 d;X��Jd�D 2}�N�UC���tfb�՝ł�31�w�8Hm�>��B��m�DnR
�r����6q�!4�� ��{�D\ٟr}x��oY�W+�{v�;:ۤXd�-�t���7[ܩX����)@G���)������B����5��u���aݺ��~�@�ኹ�nK�A*VKL��/^�T���
�U���Ge��"~g:{�\Ń>(`��H`��
����˭c=���e?�+�d�e2)���5Qqd߸f��X`�x�}NR�Ɍ���g��v�^3{������'𽺔��#�2��`�������݇�R�L���\�f��if`Y2��DQ���� �x�9�p��30���=�i���l�A#8��J�$�F�X섢�t��>I�B���le�&���t/� �Z
3DQS�{��;A�������v,�2�F��+�{`40�B��T�P��A�H�Na�&v��~�>s㵘?���6LMUq�w~�_<�(�$�A��Jl��4T}E��EM%�3wG�,��l�^7<�����`�+��zq���w��ͷ�=�3����s��u�f���1��? 'w̟�l�g�>�>����V`�晾>�W��V�o붨X��-� }�%����ذk��H�O�=�k3q����b��N}�@ƴ��؆=����Zjыz���#�6�����>���.qo�C���`�28�W��~�����il��l���PQ����R/\O�z��0��'�8,�u���� >�|��i�^ŉ�����Ym��T�d�lm��G���%T�ψ�&]l�8@���8M��!=h)�y��8�iۧ�hx�����6��C�g��� ��T��o������~��/��e*B��ݿ�����I���0.<�`E����(w�?~l�țg a�Ȕ�0�¢��z���PtŇ>�t�\�j��'iZ���Dz� >�شJf0\�R1�ŏ��utel�c:�Y�R���wDC�#h�h��O>%��<�\��t
/;p?)
�uK�o�jՐ��k�<� ��YԂL�ƥpcQ��
�[��=AP����И��E��aa����A�~� 
��՚Zv�a�̏�}f���W��[$�J�&�$�� �$ c����5Z��bq�"0����'�h�j�	``��ɤT�M���c�E�R�����a�/��[������5��1ʺ2�W��a�����ן�t&.����B�N��wc�sO	0d�nX6��{6��s_�>�'+�Rg!���\�T��-~N	@x�� H}l���T��,Tvm��I4j9t�%�NiFԀ��8�3��-xŗ͌�1��H�jQ�Z@K4�/k���:��7le��Q�N+o	2���T��@�E�@�2�k���7�������/م�h3B�����3��R������oǡ/�O����]������G?�I잜���i�Qq=Ē6���R�
R�T;�6�U��e�^Byr��m��=�dd6����0����ƽ�<����iŰp�|�n۶nk�c��s^�#X�dm���V�8ھ�/���gX��0�gX��c��Z���"~������������G�c���'�rK��8���8tA�� ���I�B&�*F�{^y�'_�{� $ts0�6�}�/lUv*�<�r	Ǟ�Jt�Y��u�?�m
����X?0
?�U ���JCJ��ݒ�NP�5P#p�Uh�sJ���h>���}t��[?��7���/��]�՟D���7a��߁b��x&A�|�@*�F��C��Бq�U����ж�h�1���kQ
Xَf���[������G��Ǎy7.;nm�x!Zԭ� ��ѯ����Ca{\����)���d����?��my7Z���C���U����\�_�JJ�4V����������Y��k�p��="ΤS, KC�Z�I�O��d2�z)��6���^+�6F������T�(ׄz��cO஻�sDJ�,��UE9�|� �� �O�S:;��cdth����ṥ�/9ٸq�LC\�t��ꢳ�m���&�F&#z$9�Xr�/^(��>lW)�)��A�\ҟ��yꩧ�찓��mR{Bk�:�:�(�X�B����O?-�)ک�r8`�~���n
�}<��}3���xD��Z� @�0��+_y2<�.���48���e��"��J�!�R�j��0[W9�'�x�y���_�_��W?����g��}�T]$��۶߸��FL2-H)���#]�\s"@�6��f!B��*����g���F~���=�Qi^��G�N�^QC���(ӊ�N4%��M�-&�����{ժ�sN���h��K�W�	=�t����L4W�o\����X�������c�ދ���rz6�V
�N!�����0��N����:�\vх��?!��
�r�7�z�F�E���xB�/�7�@��x�4|ח@V�#��ǉ��G���׼�8�;�&r�u�c����c��1���c`���MapfH�����G��zi��ч��)�?�7���L��_o���_ﭦ�4��+��G$�?~������MCS���M�6QCE��r:R,bn���/�As,t��s�0�7o[���f������c�Ѿ�+�l���mz&�-)�l�����0�,Z�ً��������`5��<��lD���kЬ��JYDк��v^���GR�թ3��o f;���eP+���W�O]z��#W��V�y�ci<�i;��?���`f`%3�(Ȧ�e@�P���+c��q�g��C^&.A�?���p�{��9�Ͳa�t�	~�Z��cbx o��,\x����,�Hia���o���?S�p�	���ox%�6��vOD����̘3�Vc��{W������6��n��Cge�-y?�E�}��M��vv&�L�$��:Ð3��k���uIM�dʭ�Ao57�3��G���w�m۶D���t�J��H&9���k_�:n��7%�����dNܩ�ժJ�}���m)O� �Z.al|D
�V�7�
|�jw���|Xin�u)F[��X����ŝʫ�	LS��t�b��P�A��;w��r_L�-�K&����&0::.	n��)Z����@O��ɼ�|�����MMਣ���F���)�c�=�t�bH]�NJw^Y{:8�9��SQ�Ue��es��Y�_+x���
�t�j�j���5�l$�)�|)zz��Y됕��U��9���?�]�;v�D�ZGW�<�����= 4S
�42�mHs��@�.t�F1w�h� ��[��k�=S�k�h��*Ȧ��>�t�N�
��+���Np��ECy����5��b�n���Z���[�N��`�J�E�L�n��]�ne��2]�z���އ�!�m�`QHN�	?w	�dx�E�.N\je,[8���c������/�c���!_0��D>G-��Y�樀�REl�9�6��    IDATB_ H>�å�\����db�i���Op۝�c�J�𩸅����ۮ��"�g��Œ�7��8�v�#Y�g��?wOO���
��������z槏��\���#��ٖo:����������u��07���ÖbE���L�X'Х�Jڰۻq�%7���Xqj �j98�#��s�:l\���"��@���j��!��kᲗ@ə�'�5<�}�b>y�f�xj*�/�� :ժ�
#�ʖ�Sr�I�H��ZQ=�9���{�����XtG:���j��"'���-;��_<�_��)t�^�\�
�NB�c�ٶhHP���+���L��*���p�g���"�Ճ�j	�0w����F�y�N�է�+/?�|��h�6��>�g��.��-Ǉ�����5��|_?�au�fԂ����FD�P:��T�LF��1M�k�<锉��8��|�O��;�i��Ȥ�;�*](&B�R\zR�,�H�!��Ha�]7���ʽ?�3g�U��sϮ��5�c�^{cނ�8��1�|�ӟS"��\��AM�4#P ��L�-���^�R1���	��|',V8�B����W �c� ��?�JO��R)��e+SיQE{{�Z�2Gd���r]�}8��g���d�"���Q�o�!�#�������RE 	E�O>��l�5Y9��e�t�"����;A^NI^��LjZ�U~PCGGN:��)&0��6 ��)�Z�|t�4/-z��3�rΤx��3f�b�%�A����щ��m�$�)��Qy�]��E��9��I���Gd%���B�B[�Co&���Q�Ej�O��0ܑ���W⍧�Ү>$�2�zND�g�a��l2#��z�93��0�q:u\t"�PY�F��9�c�I�@�m25ݒ�L�3Bh!�5��� 2=�<�Lm�m�3�����n9���Ad0��O��+�	��LA��ۿ�-̟=�c#�$��eðC�i:�UQ���B\������:& �m��1F�;��%����ўƇ�������N�2oH�,,�3[�y܎O����[�tV��z~7�f���NB�.%�W�/]��8�Kwj�u�+�?�wl��r�54�-l*���o@�pe�sBPw1#���G�C�ڈ7bj�z�~$�<n@K������M���ɑ�Q�a1�.��o���ڷ1�(�^m��w�ډ���Q$�*�/�_�u�L��In�6ܦ���zhn��~��0]�ޡ�d�@W"����y�y8h�Yp+��`��rBk��9�Evfw��i\wӗ�ꚍ���$��(�s�J9(��3�Ʒ��X{~�U�>~|>��[���mmȕ�0m�F�e�"��`�se��_��](Mb��.�ّR���}�5xA��+��_��	ҿ���.�}����A���Fò11�:�T�J6C�����Q$���k߇�{͒,��~��Ŀ�L��T�.�;�,iN�:�afq'Y
��G!�2:S�{�A���/��|��1��_�nva��y�����_��z��"��D�s��f�<99�:ݥ����e�̔n�/R�����N�x��B��T�E�����GE"�T���K
�_��£�R3�B�I���SA~-�7ׄ@��	�7l����]{�o855)�����Ь�Ay��0>6�}��W��֭��m;xꩧ�y��]BE;�ð���(����_���b��=�N7/%��@>M��<-|^y ��:�xr����v��/Nw�gN�%W��0�g#
�mk�~�+��N�&�|���0��G��C�sK"���G��G��PB�@� D4 �=���y%IAO�:&���'��w���{ JC}h�\�*�H�c�z!
���D,-nX�'��F��iJ0���ҵ�[��%Y��+�$�P��
#$ qE��ǅ������1PP4+&9�L'j�^\��;0�c�̢�h�~�l!�p���,!�|$�L
�Ø7o>���t�|�SB/�>:aTh�0���P�T*#��s��=�ɋ@��%)M{>D_��m��B]O"t�"E�m)XAC(X��t���g���P݆d����]�^���m�s���V�s,��Q���@_�/�����v���ú]9D�����8QG.���.@{���-H�,L>�X���в/�}|pudjUh^i[ã܇��A��$	�D����d\��C���} ���g1\g��_�,q��Oeoihp��*2��N��,7#=B*a�4��{�;�t^�mM�F�֭��{�Ñ��s^���f�1����������[$;�"����f�%P����Kf��~�X
����G���_��,�LƧ&a��ҩ��5f�R�Xȹq����w�6>���W���]~]�v���*N?�X|��7�8RA�v�q������Ԫ��0�ϋ%�*���V)�3��[�#�����ha�t����q��oF��eȗ}�t��:ʜv��>l��+���3��4�%�:�����~�^���1<�[��6����ի124��_��XN&P=�3�l�r9?���%#C�x]O��P� �ZY�ӲUe�v�)'�{Ӧ>��(YW���b���h�	|��G��& ����VU��$�y�-�)�*5=�O<Q��o߱mϴ���X�-�i��&����J���7�Y>^X@>��3B[�d/��[�N�ɡ���:��٢[�H�Z�Z���T�N0�lXPJF����W���ک\QրRjgjUw��E��R,��Y|���t���*�1CD��b�]\�'f����4��[�ạ�%�tܐa|4�N�8��k�]I;_���y<�1���(���s,���5pǷ�0�	�:b1�j�l�������l
n�
�M)�ݦ똋b~
�Ȕ�	��
��}�I�閭��`(a(�Jn�䥈kp$��bz��0lX�ݨ%zq�w~���7Ջ���W�	�f�0-G�T.���5	"�j	��>�}V{ wM"p]tf�E������ɗ�CW�):�t�tͥ�xYO\��������0Qd��Or�x����E��
����2m,�7�q"��jC�߅���c?t���G+���o��7��l���襰�l�
�� t�1�,��<��;��RR�끏XP�����"�nC�u�D:��k7<D�θ���^�B����g#˨��)�t��}^� *B܎�0U@*�A�^A��`�2�7lԢ��l�|���7��b���������bHW�jӚ�X*���4r�!�d��U���3QcǞYN7��-<�У8��Cp�E磭=���Mc%���^�Ǐ�C<�f ����ކ}�dq���~���n:xj�\{��m�̎ND��dv�xv=�;�t��O\�\qơZ�x9��jp�]��s_��}?b�$.��\\z�i�K�;�_����A,#�:�aH��Z*�2��RLޮ�����MŲ�z�ʦ������ވzG�ΌS�O�$t5�i,�X���
ϾZ�I
��o�Sc;0>���1�̙3�tZtp��T,�P+2��Ō���xg'�R,!?5��Z��PT)�){\��'�Y�� (����4�嘥�c���{��2y��g�"o5	hx���Ae���"0a�L��য়~� Ö��d;3##�*�!fΜ)Bn�Ԁ�X	HbjF��d�{zfʿmذA^��G+�P��u]�}|���si��[�Yj���G)��ڵkQ,T�s_h\�p)����љ��-����$��d���Ʉ��n��. �S�z�"���; ��\��Z����p #&�
)K�#�Z�[S&���@D�0�
��|��1s�|���3q��v��X��L$�u��@ͣ���j �^��L
���"�j�SG�RE!��,�<.�]Ph�˙LFU��c����fNhD�u��Ă�\+@��(:��Ço��$���1�Gb�k  �Ӵd��TĂ�p��&�K��ϲE8��8��c$�3"E�R���Z'/6#%��iG�k�R�bld����%ĺf"_�6(d؇�g���E[���1"Gz^s�*t�C����D� ��>���+0@�nO���O���7G�B�IQPM �<�	�wN�@��0B̴a�E,��ă�b�3���4-��f��qpʹ��9�L>�Qq
Tmw��m�-�0ێa|����L��5:�,�]�5����g�Hk'[���ֳ�/"�fV����OƄ#��ja�^�n�u�+p`����*�x�5���Ob|� ��3NZ���z'�i{e���SQt��O������ύ�2���p\��K�ݞ��YIm�E_��N|�{?�+��_�Fx�i����?�*N�O��o)GKf���?�����3���Oo:�e{>���k�Ig�#�:B�]M��p��R��!����R@w��O�-̙�¢lL{t�dt���B��	�J6����.+Z������L�H�"��4"x���$���W5H�QN@Ha�t��w��Ps6B�[4_:��DL:ܾ�J�OR�؝�CwHY��\S&�OL� iiZS�ZP©u'�dp�~ֲ�U�T�n���x!��SO=U		@�6mhR�l$qmd��D�>�z��8����e�y|��h���߷l�*�_�b|�C���ٽk۶m',
˩��\MiH+|�k�B�\���D^ 1���[�'�P�x�	���"����S���L;w��`�tV�ZZ�<;N��@�\:s�fR��j'|�j{�#먔�
4�(B�x�wjԊ��l���r<�Ց˻�@~5�B�$Y9��D�SW�Z&I�^9�b�����j���~XpZG'=I���I�Ha⃟&�RA  ��I~��ʌ ���fqDN�Z����s�c������o%���h�H? A �F���4�u8��Shx�4z�:�Z����ɓif�h3t�l�i��I*����a�δ���[�.!�:�p�t�����m�X���qΫN@��߅v'�ч(+����
L����
L�<��k6���X��/���`8�X�%v��u��6V�x5@��!N���(uXX�b6���>�L��}ٸ	#�!ǝ���{CK���2�#�q (#�A�B�y�7�G��^7mLNV0g�R��c��c��F/�V1^41Z�Mo�p�YT�b�
eҰ�}�G'�f��	a�T⹁zɴ����v���I^���'�=s.*��z���s��b���$��.z��o�"K@�[.��|\�{p�ŧ��6���=����~$�h��=���$!71:R]�Ƴ�K��!��������}>��G?CgWw��8zaϞ�ov��^�욨�4I�&݆�A,@��Y�<x�Oh���f*�����(Z�q;�d`�겲$�" an
�?B�H���+�;56zCR�;�����v^�U ���ɬ6�u��L�QV�Y�=s_j�2*�$ZS�A�J4ͮ��1��[&�c�#m�.���E N
CICiU�7�hK��3�6ݯ8���'�qq����j��m����P&#������ Ha��T*��[��s�=�l��J���*�������df��c!@k��z�[2::�zM�s�IA�B[.��"�
�6�)�Kj��̐�hg��H!K�Ql�|q�e�&8��̢�mI'M� ��"�L�0���b��I�����������Yѿt� a���",��%�p�k���Y	d�
�z��C*C�a�4�2�r��X��!�v�n�.6�FR����S_A�yLZC�[JD��(���9�H��S��Q\N�d�p��Lvb�f��_�	��([mh����5�+!tˑ��!D� 8�5�XyK��d1ے����׸eْ�.��M ðG����>P���8�Rf�G,�b{�M��)��&��+cz�%��"�hÚ5k�5u�A8��W��r���љ�q����?�����ۚ^�����y��������W`���Q�R�f����x�&r#�k(��Y6�J�N��p����Aze
m�.t�Xg�>�0�\�Z|�_�~��zϝB{J�����5)>�-���K^�a�p���m��*bh��j�Wq)��=���h���:���/ff�D���eP��.}>�����6o�]��.�zzst��a漽�shm�,⺇�]v������ɨT�a��9���p[�ś���$"��?|�~ު? ��Z�y� ~��oŪ4�܆�!�2?�:�Z�J�ثi��Ո���U�����G���й⎎�}�����Ԅd���������+��풅´{�ސ�@s��	L���t���K���r�.�߈�3߀�� #!I�BCa!E�F�H#D,a�^) ݞ޻�<s�ኍp:�.0'	�t���*��S)L�0�s����TnI:���zNV�|5��v�dB�a!ǔ��Y���1e�L����q��(ي��F7�/
0�-A��G�(��6�Zi�&5�V��O�3sdӦMؕ����a�|�B�6m�ƍ�q2�͊(9����K��5k�����i���Y�p������&�3\��V��M���[�\�ysg��#OI�|_�f���K���͉;�]�(�E,��x��jE
ڡ��0��P��NfP�{��k����<�6�"��i���F���yv��}H�c�c�8D� �D��N�<��f�pٹ�aŒN����*B�L�õ�$��@M���n@���pD�D<�&�!�.����*e�W�(z�tt����"J���`�X0k����`�l�N�c�<|��;p��A=�Q1�MN��_ܾ��h���Ԋ�Q�Z�+��} eLJn��[�
�_y}S��t�5���TED���Vؤ��8d��ns��;M݉�`��yh��HFM�Nb~o���Ӱ�;�2����o߿�g����n��W�x�o���0��_+�����\w"@9�P	tL���эظ���n5��ZY¨vh8v�6�0��Sh�\�nɸ�ж���#1o�
���q}alS�.]�2�lց�0�۾�?�B��V��8(�|��=��w�bxʇ���b#�Fl��O�Pj�M.�޴mu6[��,T��$��4!�m0���<�}�\�ӎ�G�6:-����w����˷܎s� _"�)aFg
�K��?��{��v�?b
���m����ފM뷡k��Q�S�?
���{>�6��G�fv��ϫ-�>���_�A���Զ�j�a*����~����_?�gW�G{[7�z?��+8y��Jm�~~ߣx������ �J�I�T='&i��ᗱ|�,�{�-X��yz[>:�7`�Ȃ3)B���y� V<��5	&�<�t\�ݤd��H�ֳ��ަ�� 9,B{���O�>K/�P�\Bܶ��+"�[�PhHb�����,��W3:(���X���R��tFO��͉���|����Ԃ ��`+��S�6��C��-	iR,��1�"�DB�~� }�ӋZ�"�[�V1g���~q"�I�=��>�����]�,�2��[��B�`q{tB�d�Z�F�&A���w�ȕ��|��"��(gJ�M ¼��9��8�5q4Y�̭�x�e� Qa��8��BS�HNi�j�2��� 7(�tJ�M�]X�#kxX��\�~�A@-�}�Z�Y��(���Ӷ��C(}��������r���:�v��\g)��	�T�]���^�H�96߫�V*
��J��T��f`����C��w~����k>\�2h�)��Q�ε�;J $)T����%DM]'$�WtL��tv6O8�m�?�Xk!bYi�#�TA��g�
��/��P��U�!.���d�|�)�6��j�E�{���ªO�'c�L�P__��{�Z���%t��w��_���DE�G7<�]�fc�������ҝ�2�ar^�WAg������Ѕ$�#h�J@i��'��%��w�~Hṫ����1������8��̈jh������<�hȌ    IDAT-�G{Vu��x�f!�6w���❋0Z
a뷎���ĺV�7���-^wCx����,Z�9g�=fZ�������?O{f��h��y�Y����\�q�)�2UE�{F3|� [���ם���|+f-m�Ȯh�̹�_�����>��Y0I:N�ĵ�\��_��{���޳��_}^�MF���>=����z��/}!tv�«���J������}��}�Q���;�}�:df.�v�S슗�0��âȫ�T��Ӂ���ft�X����n��z�p���#�2�`!�"C�"�H��V�D1s��� ����]ݖ�/���Vȑ+ic����9�<$l��B��DS`L-G[G���Ã�3�	۳m�]����?��(`Q���  Qi\���F�I��y�p俷2Vda�\�(N���p�������0-rI"%kllBvArSd�Ӑ�A'7���pn���r��B��>�m��E�1���7���-�3T�^��)ϗ��֭}��y��c�Q�\LN�KR7�k҇�W�0�9�37lɹfr=�'�������A�?�`:�V�ZQ$ay�4B�##DG�@il7^���h.�>����ر{ �>����%�F"�Px� ?�K�?�`rn�P~�\�i9�	x��\�89��A��<��v�R(���n���fΞ;�E�`�A�]K���	E�" �d�����dz��Ꜯձh��p����~[w���TZ'�b[���w��B��d��tue��5g�
M*��� <r�B-U��/c�ICr-X$@�٧�7��l���,,��	�:���������Lz񿹦�az^z+0}�������+�q��h�P Rc���Ω:~��:��6��Z����e����Q�܌�9j9��a$���j�w0����.P ęs�_|�r[#j1�e�e�H$tdg�0ԷO=�"���e&�[���-4��c�Q	2���L�1l�>�0����ǯ�cv�i�+<tj����_��|v�J|�[���NM�4V�����Ƕ�Eo����,�P���[M�n�>������'��g��6P,F2Y��yct�]�B��{F°�O|�\����d�Ƈ�(б�W�:�����7{�sF�Q���\�q��ǝm�@���n#f8����\�,�����^{E�q� 
Lm��Rca��XY+MM��u�X<�eo>���������g�G��	�Ђ�-$ ��[�eD0��ZЛ�R|�2mi�5Dg���=�p����k�ϛ�Qi- R+��!����P�4�&�G��P��Ԛ� U��4'jҐ�bS�j*�\�(���T�i�U�w�F���5)���V�����Ԁ�.�૦�o+M� �BsR��n�BiE�a�N1'��r�R��@',-���^q	Cd1�r��X��� ����4,N?�����1�Z�� H�3Oޯ�/���S��d��Ktl2�l�`OÊ��2�jD��/W�qU� H3���N�5�O,Щ�B�.c�հ�� K;���lF����̓��-�}[���OE�֭Ea�FW@�S��µ���	�CQ�6��ի�4�L�e�����ׯ]�3��裿Ea�C�=X2�մDR��@�Q����/X�b?��f�x�[�p�Bn�y�;p���๵[q�eoCd�K��\�g�Y뵆P��'D��Bq�Jp=%Rދ������	@����O8�\�`���]�V&e]�����`��N�2�������?�_į��MO��Kb�o���i��ɿ�
lذC���[�:\�/�،�6��0�E����5�ŕ%c�H�9�}�J,L�pʻ��rHhU��e1�l�F��e��� h]+���nb����a��	;mb�Ƨпy#��E�eڥX���rPMl�9�m��P����v�f;�
�4�%W]�ם�V�Ez�*NU'^�Xܚ;� |�KWc��������U���F����ś	��
�+
��5��է���ނCg)�y�]z�{��o;�����D��⃗�RRS��P�c���h��L�j]'����~|��#�h���P�*���L��5~?���H���wGo������bq���(�V<���g���R	}讏#���䳲?g��cя|2ݳ���p�Y�1������9;�I�1}]	�ə7XF��b#��@TW\:���%��1w�L�a�P)�Q/愪��ǚz[
e�n�	m�|���8�ҭoNŊ�VS��+���˖�\�(;a���A�Hm�|~�J����W�kU�Jȟ��$De���=Z���J^W�"]y��B/jQ��?���Xi��S��
͉�uCC*����\9{&-�R�o���r;P���z�]{0*��A+D�\�?��Xqɹ�ts�b|GȜ��~��!�T׆ X$B�T����%.�I���9*AXҞ0��\�~��r]������!E�H�S �A�_��nj>���&V.ݥ� 3���5-�IUK�c��!��ӓ�~P� ���9���E�}&��Sǭ�p@,������BؤJ	4����j@,�WE2n"������QG�-[��]W\�|͇�"�m�SYxuW�ON8ux �,�y�Z V�&�L�j����|UkB6o����k�"�8b7~��� b��H��>|z��n�~����
��e�>��P+�~��(_��痳���7��X�}~�X���B�gG2�VQ��ȅU�����!�0'��(���#�H�UJ��Nc�A[�LD��Dg���J��w���p24�L���7����t�a3�!v;wlB��ub���h�N�����j};�0V���h��	��+Sez����P7��H.CӅG
LV�ZӲ�Ő �J��k��mmt��Pu��޿V���F�N�	���H%c��EԽ���1���}ѿ��r2m�hD��J��vC7|\�����#��.,n���ϫm�A�f�f|��e�X��L���@݅��ƖT(����5_�K��J@3-.Gr<D{��u�{o��Ru�U\x����3~��c�Μ�z���8 ��y*�u�JM?$\ F@��N���	��CTn�R�7`H��BR�Y�6]���60A/t�����C)�CX+I^B��R�3PR�O9>����#Mg#E��s��<�]x��o9 X���\W5�PT�kK$̟[���Zz�D�cIy>Y��Ĭf`����o�Ⓒ��jGT�]U=����,$YL���ajB �h��M��(U4_����M�)�! N �=JMlZ�V�3�8C��;;z�&�����GP3K�>  ڐ�AR��m+P�a�&B�9�*&���)Xh���� ��)ݽH�BļS��4x�ݕ���v	�<�x�&G0U���Ę�#�[\G;�@�^���%���u����lZ?+#^?�u�;
��08��5�ʚO��+�1c�rl޶��Y�\�>?]�	���Y,�����#�O��h�`�ޭ� 30o^'���K��w�L��J`ϪɝO�K��:ˢ���
�ŉ�.d=F�-�UW@ݚ��x�̙3�aa�����7m�m����a��!^q��t�0��
L��t�_��}}���R	���А�z���T�(Vo�X�G���BE��p�F���7�Хݒ���(���Йf����bђ�h��η��3юT�L��䗾�Q�*ŗ*B��v�����(-O�\�cp�  .�C~��J5D���Z��C���=��P�:)�]`h��j`�� ��e\�����?��A�P7�/���R֖NabpH�ot;�Vi,(�L�U:���h�z*���v� �o`����'>4��Y�c�'���Anj�}fq��{����цl"�b���Ys0c�,u�yu��h����	��	�m����IS�l��
�$�S$3$���<^�@Q{<v�+e詤�3 �5���# ���R�	�+�a�;�Yq�~->��g`;���,��}�	�Ë���)�mФ��Z
���Jb7������!�/�̂i�h�u���&��5�mC
E&B�N��7L)�Ӣ� Fw��/��R�)�Q+��;-���xk���%�� ׎��[���U E�
�J�l*�C "��;�I�X��g9�L�m)�5�6�iF+���&CQ�4��(��
n���~� MM��Oj*�S�r?X�Դ�h[��G�R�	�a��SO� �e���%oy�Y�^���'DS���FC��K$�0SI8ts�u@��S�MzV�ё�)��=�΂�3I<Dd����4�|�[񪓎����ƇE���EH퉻��P*��D����b=ݚb�d�H�9q�q*E ��e� t�i�F<����u�c9�OV�윋��"��.�@�4��nNԗ���1���Zb\P�A{2����L'�;����o��[oG��Հ:N##��VE���9]&!�լr$ZE�q�j�p�R�&��f�M��E��z�����Mt���ò�m0�S�B'�t�Y	L��b�o���*O��Kf�l�����u���a0��C�<���T�@���/M):b�ZuR�i�9/��I$�Id�*R��ȤhkK)ZH<	�c&�f͑B��yR�����F�z��&����	)4��"�1[h&�2��q���*>vM��3_A	D�.�\���Te��|�O�>�*�$��+�"�����~:��]�&�T(ˀ\pe�$�L~�{���O�����k��vkX1�]�@��/�D����A��ŨƯBo��Q��E*|�2Xs� �Z��b���݋��Co�R9 �6�|��C���п��s�(DL�Q/r"�P4
{}��8LqzA���{J85,|Md�IT�9�'�F��J� �2��_�)mq�OB��FUǕ��?|S�vq%!�\��%��׫�0#t���7���^ƯQ+�`�.b��l:-Z�ҍ�y��ж��f*@OM.Z�kRq<Z��
P(ʒdY4�P-�(�`4�B��C�R�
nG�<䧊>��E�j�=���`Z`�R�0�k��& - A B�5��:r/�2S�H{B)��.��ӭ0ᦛiX��PʘH�f�&����\ �A��N���ӫ��kp�ði���� ~�G�i2��]Q��x��Dt�RŲE�ёƎ-���`t&v�0#:P�5Z8��7��y��8��Q)�Pw+�.Z
��P�ck���s���:JX��-��C�����ǎ�^���ZU�^�,�|�9���0���wѾ�=�>Gri����d��3k0L�RS���{�>�t	�r����~�˒J�Ϻ���C|�?E,݉��=F0Ͷ�����_lu�8����E� �iσe�8�&`L�n����P���l��S ���A�Ґ�#��M�b���@���SN8~��z�|�O����
L�<ogdz�GW���h���t�B˂���1ZŃ�l��Ƨd�"�J/y~�
����f�E�)�7�����a�Gѕ�j�ϟM&��Kqz�{�f���(Uʨ�H��2��Z�J�0��e�]qf_�:�Nd�\G��)�����k7c��#t�0��o����a�L�P�({�L"_Y��Rમ*�Ia����m�a6;�:���[��y�����nZj���f�XK�����qS�@;Y�y��ɴëyH81��Q�I����"cI,��j�6#?�R� � ;��O;a�m��8�$L'w�;�;ԛ\�j>L�	�1bI�Guݡ���A `��Q��0M�6j��J��Lff�5j ��48ٌ�^��:�|��=*�+�>E�jf�0�M�M�� ��b��4	|ޒ��>�����'����Sm�ue�J0Ɖ 5=�_�  �YD�8�h��G�� ��[�Zṩ�+R���k9SI7Y�t�ʴ��.�B�\��%�ѶAq7��	Dc���ӂUB�te�+4�f��l��
�00�E�b�F˭���5�A��׀�H����0��t�._��*�:'������s�A�#��
 �<�`���r�妊x��Į�1��s�E0.�MΣ��w ���H�J���b�=�$9˫�[]�]�{�l��Q�B	�E�g����o�>l�`0`cdFB���6H�$@	P@ $��Zi���qvf'v������V͎|��8����lOw�[��s�\��jhИ�Ú��q`�ԏL�L�X;d@i(*!� Ǯ]�?���i��vkN4�Cc�͵��TJ�8���4��aB�dNSt};6�V[�)��`�R�2���(�Zھm+n��v�;��A����U�s�8�a�Ie4��,2Œ�N]^�lIcC�N��'��9,[�W\�,�G�:�/嫸����?*����Q��8xP4;�E�3"tR��df���W˜.0 _�4�!���>�E7��W�(�&k�������ї�����'�]ǟ��x�y�	ȯ������
� �S���6����v�v�;���/��"6m?�;7���#m���I=�5�6�>S�מv�����R�o\�P0��N� r�4*i%�B�"�;�f���ŋp̪��:���
��vB����rf!Ņ��]��s���i'��[�t=���i<�{���n�Vnv~�v/��14.�f�΍�
L�5n����l?*�ȗ�&��h��W�Z�^k`�6�\�.J���?�	מ��,r(�5 �8��t
b=b�`D�djM*�lى��)�<����Ib!�"�:��
b�iCq�-a5�J~���(&,�$��|m?�U;h����hMM�����U���ϡ�l����i4�a���PE�s��P|w"R��� E.!=�o
�F�Le�zQF�	SB#�h6��9�����������榱r�d�!\'@uv��	X��"򙢶�oQk64슬H���Ӣ��ɤro�;����>~��dAO`���;�v�Ʀv�:g���~��?݄h:��z�) ��y�k#W*+�1��k���k5y��C��ͯ����U�G����D�Az ������ۗΘ�"���������\'b}����Fv,��y�C@,��Z�.JeR�B<��q��/��w�	�;��~�ON�Ns��s�[O{����U,���IАgi\�$R��%�l�Uk0y�&���� ?
�HE>���qkW��o��nX��w*�����Zw�')K������i�֎�#���L�hNx�K��f6��A�Lkc�K�|�M������8���\��)C�ix��Ӵ����C]/H4��ũO ���.����*�Ϧ������1k�"�,^��E�x|�V��F���_L�@Y%]:�J`b�����~F�r����D6�0B.�b���H[)<�iʹ4��6^����K��VQH[8�̞������
� ��α���ϱ;w����B�����i��}xt�f��N`&
� "ߟ�A�)��D)gaq��i�.�p.@>��ۙ��>W��)�vͩ@(�ɉ6���b�t�(��g���Ȧ`�N�2vr���9�g�f<Nq�~U��l��C�N6��]C��׼���Q��� �}e�f)��}�>�d'1��,�d��b��k�Y^��Q*�M�0\,# ���Cw &��E.iO|��&0�Xd&���,fR���d����2�- =N��f��B3��#����Q��$j�G�v��s��-����ns6�CkfFx!S,
����|	��-�@���-�ȅl��,�m��v�Λ"��ҡ����f2�М��Ju6Bh�tò��}i�v�h5R�.(xHEm�M�C�N��8`R��2c�=B�������,�I��###
Lǅ�Ѱ=�X�'!J�2�"�mµWBv�$ "�Y�A!�7Z��с0�;����f,^gFI����q��z;i�L:�@D��r�"�,��o�l���Q�n����0��O{^n�Ҵ)�v���!������g��]�A6�G$�f^��=�M��bQ�ƛ��<��O��K    IDAT�-�+�/�0��n�QZ 0�2nc�	L��e�b6� �v@bJ�	lZ��8y�Fԧ��{�6�:������בϤ�r�(���ގ��_���VYڶ�5%�'}MH�;��jy8��ufl�=3���5���� ���P	���݋���z>�0�_Z��:�wN< ���!����;�%�h�t�CY8�:��:.{�;��C9��q3�m�15��볹��%�1R�r�,(E��2k{!�ic1���&A�����[��1���w��%�8����k�#�l|+J�����7����c����Q��8�i��j����{Io~�
�.��y�[�+�c�hlb:hvBt�yl�?��؉��0��,�鎤��$s�OZ�j� N*DmlX�K��v��&q�1��u�M�G�	Q!%�beY�23�#R@��錴
,��LV�;�N͠���*v��L��"�l3��z�C��E+p066�F�]k3=�vآ�D�@p+�|O���'��n�l��Eױ���B�J%��:��I�6��t�ظ����c*���`7�I�.�,-o��	��V�]�$46` �)�j%JL�Ѓ��b6��禓N1�Ѱt�ic��V���iy��g�V��Hl����H� �	Ų����1EaÒ�S��Ƶ(1��B�ΐ;`��"�L�&��o*\:�F�	��I���i뜀&\"�3��
�cƈ4k�Ck�+��������&��݂�ɉ&��g�+��l�Ux��N�h��0�Dxn\�\ٯ�8%:�{1_P�??	� ��$�P�w�:����Wtv��~�3�y3S���X�x������*�)
N�a��8�ä�gE�"�n�Ȅ��th��I�8)#h��.Z��$�� y��C��gJ+�1hw�o�>���E�ᶯ[�^��m�fsX�j�y�5�-,[�Ͻ�"ME8}���/���A���Ԅ�1��o^N�N)��S*8����d#�;i��'mؠ	�c=4?1�0J+҈��lxW._��|�1ܟǍ��:���~�J��y�$���]��<Gyǖ1�&���ł�$?���h�t��.z�7oy���?Y�b�O!��h���@� ��"�ϣ�&�k�B��Me�lڋS������߾�9�i��MG�BQ:�Z�-+`6�x�	����ߤ�s
�V���G5:��T�:�?yp.��_�u�6����QO�],:�.vl݊b��`1�?�����K�t����x�٧�j�^�[�_pz�/�p�_��\�]�DO"Hu�B8�>M@�y��ҀpB B���}��m3e�5#I@�peRz��b���1#9d<���j�ß=����|�c�����tZp3)�w6�p(l�H=ʠ��Z,1Ұ�&f��}�ƫ>B��tq G�D瓵��:��n"
D��Ts�֗����,trE ���舴(M�|Hg^���!�I�}O�,�Oj(1��h<�Ǫ0�~��c���+�O-J#�V�X�?�hH����E��F�/m���OP�
K(N��v�� ��њ��R�� -Q��(��vŅy�B^�ԝ�֪?d0|�ԃ6ZՆq�y��G')&-�3�N8Amvc�������0�J7�}'�>��6�0D�B~�\�d-���F.�ȡ}h��`ώ�趩�0Z���iLL���a�������v�Z��ػw��j�����z=in*T)?�m]t��'	��߿�w�&&�x�� �_���_@���,ho��M���t	X�EZO��U���{��$�4����ەA�"K�n�����V�^�����x�G������������o��zm����җ�g�u�l�"�;�߿�ԛ����矏m�?����:��+8�� ��w�w�Z�d�����k�	]��h\���alyb.���88~�6�uc�eQN�R��
eQ=;�JJkC b�Ky��6t��nB��#?���&�[˜���m��ڵ+�?�i�x��b�a�p�FMB8���ϥ1��Is��08Ч����������'��5f\�� ��_�F�zU���3����`ǎ]����F]�3H9�w��:i��&����8�E�"}�-��ЁW���J����8v�R�I�L�8�*�&Q���ca6+O�Yi��]�9)�˜�T`�a���Cd�R��M���|�k�s�0R��rZh�� ®b�m�;�J.��W�k� �O�`�x�y� ���J��W����_�*�>�)������-���� ȴ����y'�~M+-H���%�����i��Φ� �ʈB�M�6K6F�6���(��(;lN $��5�G�:s���A�,�S�ap]Z��~dcbv�v��Ek�|�mԼ�� �V�s>@�U'e�>b��,�,�c�U8�30��%�115�����jQ��H����p\�2FK�Ӝ$&��:'��~�K�Lt�Tq�:C�	�`�4-i�9�I�D�NWt��K�;2'��P#"-A�r���P@��b�a��6�����"*�?�qj#! ���f�J�N�k8_@��tEԫY���߆c�VҖ�Z����8���<6��ɇ�"��2f��Sq�
��ְ@��yІ�P�2�.F����WA�]��	179��CcJ��d�B�G~���d�.�<�T�*�v��p����Y�8_�o|�����(�;���0�y睏������رc�@������5���{U|�\�J�+��:��������Z���~���| ��S��R3��o���~�����^h}���Bل~�?���~;�f����
� ��s��5�^g]���=��G�����S�����;��c���K.y�q���o}�[�RK�/ý=$�7��Yg����w��x��a������71>6��d`@]��K�KH�FC�+Q<
�>|��7���Q��N�4#DW�9,i�1 ��% t��
��nl���7F�c׬A�b �S<苔���J��9�P_g�q�~���xt��dk[)��p�Z�rpV(Qo��:�|�s>��Z��91u3�82%PG�l��Y������q���ơ�)�,]![�L��\m�yfzK �uh`A+cGa�Կ��}.h1UkW.���Ь���E��Ǒj] $M׹ZYf��8�JK��s�����֥Y�h�7�s�S[���b���>�/806:���l����[��G
������Y��O^�uKa��`w[��g�D�O��{oC�V�@~�Io�~�+���}Q��kuqpjv��n_��.���Q��(�-d�Y�0���Q�N��Ψ����m�GX9Z���r��W�M�o3��J�J�� ş,XB�݈@'���bb�����E:[��u���'�`lra*���������,�3�.2|�ND�~&2�6��C�+(V�������5b�yp!J���F��BY���e����ŏ��D�%W�@�=Q��Dp�Q����s
��-��fs����p��H�fdP�ҥ}��u�V�`E���T����aMC>(B~b�Ϣ��ǵ �j|6Ҳ���N��#(�od�X�4�.�3"vMh"8nZ�^,�H�e-0��$����� �L�J�"g�X��χn˖-E�Q��܄&_��ѨN�K�CZML9�Ç�Q.U0�x<��|�2�LO������ۨ0�͏n���E�(}�kqه.�F@�#�Wt:x�ހ7��Mh�<��G?� (��+��;�St�SN;U��C�
�{�^���6�9<����!���֢��������{4ač7ވ\� ��n��>����6��g��4�����K��6��}Gt�9O�ҥ�p��P�븦��+M�.~�lr�=����~��Q����5��w� �x6o~T4�B�����]MrH�l�j�����luF�&_,��W�L�LoՌp������%\�����ׅ���rO
'�X�iX��
��@g�qڢ�IdFu;U�y>{�Z�P��#�An�F�Mah����,�m�/<����AM@Zu:�y:9A�yO��a<δ�^�h��"��.6}�G&u]eWQ}���ҕh_�k�.����w@:�O?�۪��@�n
e�c�3�H�#�+�(� �L@"9��rhuZXT��s�_�b*���!�;x ߹�N�M���L3�U�d�YM���J:������kJ�D]����)���v���Lϡ�߯d��Z]S��RV�\�{�[� ��Ji��/��c���gy5���{5ԯ�����
�.�����m�/{6o����O��J#����-��ݻǖ��h�6:,T�B���#BP�aQA�f�m&bS�M�Wڅ����]d-O./���"��_ʚl�(�����Y!�`S�m�*u���&��af���Z3� �s	ӛ��E'�+2���P����U�u��Q��G�܏Z����8t�"�#�^�u�IȒ����+z���Z4���C�e��>�Lԙ �4hME�5�"Gb��9���m�� pJG����Z]�o�� =�9=aj8��*���cڿ Bq3����t�
<x��p�yd,^���R�aeX�:�-�;�t�Y�j5��`d�d��Z�*=M���2�$|�3sѸs,69Qq3�X6����p���@Ob��u�&F>��p�������Z���)4���_p>���+qd�B��)��.TH~��_��?���������'����~�vǭ��P�ڱSG��w�[{9aQh�����Wⵯ}��裏F7�|3�8���k��
n��<b����;^x!N>�$i6n�(j�g?�9����q�
C�e����S���&�~���[��؍z�k��Uұ�h�d��u���{!V�X�k��5�u��(W���;��׾V4-��S���^�J���/�米_�5��c��G��^�����1;SEZ�MM!_@sj
o�����q:N<��-���us���݋�{����������[�|I�Z��qBB:��nu�Q�M RD*G�(�s����)o��H�x�N���>�H�y ���-ڪ��؅�Y^���5 e�'{hNmҋ^�2\p�8|xB��Z�T��m�M7��z�z3���:^G��J��j��N�ªUk039�F�it> N<� d����[@���a�Y �6�{6�<L~�Ec`f�E�ۂ?{�y���?|�t!���̗����DxA�4�3�Ы�g^9����nN�����.pfJ��$��D�;�Qa�I��d�������=N@@^��ḕ�p��M��z5�/�!�{�ߙ�]<�3����?�
<�yktd��(â1�ɺ�����=شc��E�'u'�ͨ�g˻# B{]:сHD��cZ����O8,��[�*e��ie��J�
�s��b�ё����>�wQk��..����^$��d��J�9И�!W,��A��ް���2���/���G!�U�dn�V����q�B��D��}��# �D���䋴w�#�`�,���`w��ͣ13���`aj���A���0�`�>��n��,b�W�iIjz�,�sA�}e)���&LlK�sM[Rm�;�a�m��M��u��n6��9�a���h�*f[(��n�U�#����k��պ64*6,:	8D	#�0�GO���G<��:�O�`Bz�u\z��/cfz����Bu��n��v�޾]����s������K��b�avv�{���n��6|��+�E��gD�W\q��l=�ؖ��^�N8A��×]����� :��m��(^����g��={�`ݺuY�_���g?�Y������.�+^��֖�6G���7q�i�	D|��Wi�l�M�L�(.~��q�%���O�>��ˣ�O8I ����߼�o�-�7���u��7]�������C=�R��V����u|�;ߕ�����7�ٹ*���,N���V��{�Q�E0M(�����h�	/NH�I
\�1V�Q
m�����*U. ʺ��	��ݩDK�p�#��5+W�5;�ݏ>&��rs �����:�P�g���=��F�V���\��� � �Lã#X�~�>��&<�������xl�h�=�D�5�$���%2�v�gI�EAY��FW-�i�v�8��+͠�r�谱B�v��);'!���ٌHG�s��C��UKP.8�蕟�5߹�0� �ˁc�	��i��V��*ݞwgKhX�OA8F���U��jc`��6P��u��)����K�m\�T{
~u
/���^��<X{����X����;-z+�`@OϪN 2Qm)	�������K�Ft��RE�"�\����v�����L���#�N?���(�@��4EY�e�=M��	F�`^J�h��O/�@V�z�ر)�=&��$Bv�ʦѠށ�t���u]iY� Ib ";��z�����w�:*�pQA/b<yP�(ݢX,�"z! �Ht�b 2nS�h���,
n�٪���G���1B,ٰv����x��bȸސ�FN�� |�r�!@ ��π@����h[��]�J�e[:5�ծ�e��,�ɖ/�\��i�';d���<�g&R���tl`|��A%��v>M"y��E��̳���E���s��-�A��DJ�����T.��UC����K�����u��*%L�ߍ|%�_��x�����&��S�i	�� 4�\@�������mOD�_=6w��ؗ죚P�٬^O:u�,_�?��?��u�q��A,]�T��+_�*>����$y� �կ~��s��7܀�;N��O^���w�ѐA��u�xγ������8���O\���SO]���]�z��A�
#��{׻q����ٶm*}��>q9���[�����:(��lx��u�1Вt+NĘ	C�^���Kz��D^�VW�=�r��G{̴`1��ë2̙���@)+��N�|��Mc��|LI_�|�z�}Ԙ)�V��f�L^Gr�����d��D������8#��]�(�o�U,�B1�G�X���{11v):mq
&�`CM$m��I�A�˜��8�Xf�N%�+Q7y�d�yF�  ��Q���J��2��Q�Ǫ�����?����.�0�u�O��[�zˆ�ax����@�y)Zh���]�#ՔV-57&iit�%�tP��1�ׯ	�ġ��Xr)Q�N]��?�N}_؛��
��
��+� ����~�r�l���F�$�f����#�����G����6)0"|�5-�hҧHM2�%�9q>�ڂ��ѥ=�~)�Z��)p?�`����Y�ĂoR�4�����ƵcR��7?�`A�i�K��28�j�iD��ݧ�!1�4���A���1�Z���]��37����*��'?��m<�H~�tbR�Ҵ�d2�n}�26�Z�����Դ�c!AD���.~�n�-�����bAH!������t�mt�6�u�޳0%%�tM�l�$��̂J�)���)dW���!q���Ϫ��瘝8��^Vl[\t�������M�����QΠ	�SȂ��Ʀ�.1��}���	u-�֜�� ��{�z�n����UEzx��.����n�O}"�P� ��V}�RŠB~�11�C�^��7X;�o�PN=�T�?���>f;��@'t���?�3%�����J�������GW+
�[m��G>�7��ϭ�{wG_�җ4a�{]��O�� ������Yg������������W|$:���]����я�K�xn�o31��;��ע�<8�C�a���[��f<��!TF0Wm��7"j��1�&�������X�NK�R��(=ާ���� ]0�K�ZR�x�ZȤsh�ऑ*g�ʧ:IO
P�s�o�V�\��6��E�\�.���<�y~����w'��s�������Y� ��ߤ2�G�Ц��N)�f��0�㓘;d�W��Uf�G�$ �&o�������%.<�!;
@�1Z�1�l��N#A3H�>�5K������"�����[�۷� ;�����oN<b���R��g�����La    IDATE�F��n|�b
nK�;��R���5Q?x N�E>��x��5�p�ӈ�5\��g�j���J��S���]<��U�}�Sfv8��Fu�������-?���� ����HI�m4�A��5~�Ŵ,u%��$����h%q��<��p��<ص�&+Bz���$|\L'}�q�Fe�b�+S6&gg�	�$�\$�c�@%�P|V��?�$�L7��' I�IEtܑL����!�����I�d�Z (�9�8��~�)���c�l�����^���a\�ɫ`gl�8XЋlA��-A���o�L��[Q`b���u67NL��`w\�*�t�R(-]���Q���!U�6A�ܫux��d%�C�ٌ&A&�[aolɴB'D*
��O�(��K�,�M��Q�a�3��2��:W"���Ki�ԙ'�d]��~���k�93�?|�Ÿ��/Z��ǣ��N>�d��^��Oj�)0f��m U�mo{���c=�����k���d�{���<���-zHW��=�yx�߬�5.Po4�{��w�w�|:��B�u\�/��^�zk���g>�������>'w6ҵhyKN>� ��_��|��J��>��ݏ�n�I��ǋ��}��_Éǟd}���Ft�Z�d9������_b��A/���,����q�1S2y� G*��FY����R4��>G���
̇�J2hlN����E�I�NkR" R*�.��c�%��%6@��SV� ���7�Uȶ�2�+^�l6$	�n�a,�	D��0P�[C���D����t�b��A�Î�a��,]���q�~�qr9��Sp
�/u^kf���0M#�7�ؼ�c b���=� ������S�r�*"o�����p	~����?���[F�w`�]t��ܯ�����KZ ��M�n@�1� m.D_��<Rد�ŢJo�ӗJҭ�#z������PO��{oC�V�w�������ZW`ǁ�hbj]+D�6��.�溸��{�s����A����rsҡ�,�&��P�H*�$�����۬�Q��St�R����5SҀ&�prLǞ�Pz-��,��|Ѿ,f��*J�p7�T>���EHeҨ6hԪ&X�t��}^�����J8~�lmM�e\���'�*Fg���4�1e���N�8�w�I����n��%KM�}p LǮ��r쒣	�j2c�i�t�j���@�9/���Q���	U��^��;Ȏ���xő!���e(����9�o�@40�w����P�b�>��`j5�d�Dt�2S.3����$�$�,n]@�Z0qR�9n����ʭ��08��:�d3�����,cz�^���_��u�WF�}e�t�ɲ�}�߿W�<N�� �=�����-�f��G�~�!���)���[n��'�ɒ�+v�	:('E�?��(P�Dx����?��V���E\'���q���O_�j��-��뮻�x�3�u��WË�t�c !���O;S.[��}|�v�e;82=�o|�z��9���+����ֶ�[�-[�j?�537�w��oq`�>�,�l�����Z]ԙ�m�F��k:�K�_;Q��5k�)5#�pO�	��b���H���4=R�Fp�rZ#^Gi��4�F]�~�)h���{j���}!����*1 @���{�V��5�׼�.*˗���5��TJX��T�Ʊ}�&�vZ����D��Bu�v����E���,a�X���� dp���asЬ�no4���9s8,4���W���.����v�ձP�j��l��O�i%���4@8mI�-�4�[oǎ}�}�T�r���˖)p�����������K�a� �ك(9!�qΙ������}�Syz�S���������툦fkH��B���L�ko�)?0�v��� Db�"m��Ǜ�xV�=V7K�a��O�@�E������%��,#�	�D��.������LfA�
�E۶�����a��L��@i
U=#�f�?����3������U��Ѫ$���G�ь�� �T%:X9�+ ��*�e�[��蚵*ji۪p<:�d]���p_:!X�D-�FC��ufhH��?�L;a��kz�O?ՠ-�]C�$R�.�=��S����6f�6�v�n"�T|�'ϩ�D�b�Ђ�Ǉ�Vs|�F�dʱ6��pĠ��~��wPu�- z�v͋� �����X�wE�q���൛�+fѪO�/��\���YW^yUDa��U�08<�+>q���8AH 5?��˯��������Q":���߼��,퇧��H`���������u�g�5J�8����{p��+�O�B�P�����q���+��`�"���9f%[
�C}���w���/� ��l�"��037NP4e�!6�ѽw�;wn�]x��ׇ�|�}x����+�"�.B�M��>I����&�;圀� �x\ 9��JH�G
�3��'��R?�rI	���ś���hA����y���z
��9<�c���ӘH�5A{<��y�)X�Ѕ�j���ׇ�e�0ݬ���t�5ԄLNc�}����D��#� Ib����c����$@3	Ք���\M������CPDJ���ɜ��b��#�h�Q3z*�F�!��n���Ӟ�fQL�9����?�^��1}�'3:9��y~��=�S�b6�+V �ؽc'����%Cx��^�uK�k�(��~Z/	�������
� ��̡���ϳ�<�9�6�H�����o�۷o�3hum��j�ӗ����ju��>��2]�yzQ�t�8|.	��30�N
b*���Ӆ�>@)l�U����eੇ�S�a��՘i4�h5�!Ϛ���B����ւ�r��9E�&��z�����&)�����,�V+H�h-,ү#�T��D�Ợw�~A��ӵ� ~�*
G�V�*�(T�Y
y�A�VGmr҄2W$!�C�����9�j;N�"٥��|O�����NB�k����l�~F��uD�:@��W�W� + Q[�l�ج�-Y@D=�cKp�&�h,���ib�0I��=ֆ�	��6�~�9����n��	���G�o) ��dL�{�������.�^��߷>��/F���B
˿wۭ�¿�j��
B�,�~�װxd���D�b�k�.|��7c��=̓�9��S���W 3@̿�ʺ�󟋸}�w�T����O�VuQ�l�O^uN:�$9<�,�R_Eߩ1ɰK_�`jvF���^�r\|�Ţ��?pH��׭á�c����K����4#��s�IT�T�Z������ɡ�hcpx)�jMIz$�ָI�jf�cW8�.'D��&i�HjÉ&D�b<y�) '_��g.�}���JڱQm�5�������,&��ױ���?���{�3nn����\#H}WÂ 9�j��6�@1vlI��Ԗ��uQA���AR�V�Dٲ���o<
�)�6&�qF����2���q&q��j! �dxD ���ڶ4�fL�A�絍��9>lp:�vD��zE��rE
NK5��0.}br�^�m3�� xso1b��CX^��q�*��`��52�xb�6�.��m�*�- �	��3���P?σ����
���]<�Ӣ�V�'n�m�b^����'����vb�DS9 /�G�"1L�/�#�Ɏ��fG�`R%T�����)C�b�͇!|ȡ&�tӎr�c7�&�;x�C]�ZXJ9�n*���D@6����P���ɽ�yJ��|�	 I��^��t���� D���j��|�y���p���W�>��7�)�%�(3T�����B����%L\t�����Upg��_�!��U�,ו���'��T�vF�I{��l�CX}]�^7T���,E�!����{�S���~f�9�����u���`� ���b�������yA�q�J�R���	��]��׊�1 ��lh5U��O��&~�7�~u���o�����9�dlۼ	�8d���=�>�b��@����8:�uk��}���������Ɨ��صw�lKI{���MgD���`��8���,m[^?��ݸ�{t��ͧ]1��.]"Z��� پ��������ls�o2�33x��^����%ؽo-Y���G6��w�{>��/|0e�:;��ϻ���r�����۵f;���Wc�ހ��an��%̴�i*X�L-l�ry3N�Z��(mR���Ф�@� ��u��h��H@2'$��Ң�p%��u�%��/�yeW<�׭E�v����Н�2�\���99�w��N�N>���Eݧ�+TN�x=����ʻh�*�W��,�����Ή�t�RR�$Ro�5�kO���� �ɾq\���!��"�����]yJ]X��(�5KZ)o4�F�(��$(���b�Zf��cF���:37�@p�c�I;X�z��۷mC>��p���\�:,L#ݞ�4�̳���PO�����[��z�ϿV�W����=���*^�B�����x`'��E5���U�T�c��'�% $���ul9(��u���q�uR|��bޡ���$�\b�@�]r�t���Lw�8�	��c�8�/�n��j����(�� :���a��&L��?�~�_L�HiXf�N���K�k������)����������h!�J9��z�Z�*;�t���b��x��.a0�,�V�u8قq�����3܏ʒ�F�0[�bnzN�����jHuB�Y��IAh��h�E����P���t)^�Bќ#�I�p$|��)���� �ac
_BKhz/q�H�YO�B�#+B.�,����VG�)�����XX4:�=�@��A�Dꙇ����Zv�K�Bl��̔���ع���}{�JC����[��mwݥi�@��]��3k6)��v�#�Q�+azzV��(����f��~��x�3��'�*�A̦M�4-98qH�o�6�b�1+����$3Et�2�~���D�<F<����.ϱE5�)lA���<^׋���l��g���nI[E��hKf���<M�M�#S��ֵ';ڄ��&��e+b��Ѝ��K<�2r�XI&���鴍J�(�7v�B9���h���|�.��-0n��ۡ�'k��SA �)�5�4]d� 78�f�l������o�X*���OG�I��뮃7��ˋ'�)�6R�#:$���{K�ϙ�Y*OPD�D��	�O{99	���'C&���b��E��Qgw9��Ҟ8�G#��Q����$���\��k9�iA����[�>��ʽI�un�_�F�,3Q���u+�׼}� �NQ������^�;P�v�fz��̺���)�Ԁ��k���g9ht,<�o
߿g+��F���Ǵm�S��sq�Z���#�0�x)����j6U�Q���L�����t,=<e'P�]H�WBFS��j�&Sh��ۙ�K���|!/{�(M�|�OJ�f�$p��/C�J���2�6 I�r���$ s��� ��c���ʌ�LA�/�1����t"x�:�f���$��x���F��=L��z<����r"���!&��`6vikZ�Q�	��z�ze:�=�����t�z�c�1v� �,Ӯ�/�p�8ѻ��bw"�A.��%�0N��	�S���ג+Ͽ�3� 4Ѭ�����ԦT�g�cR�M�'A�����~�J4�f�w�Nx~Y�YƽK�����v�[�:�u�M��ݳ�&"<�r�5���E�bf
k�B.��Z��ti�Q��Wם����0��S?����2\x�E��ޟJ��~�:�q�m��{����A�g�)����7�Lda���hx����dA؍��./��P��O�Ȕ�t?ܖ\6���iM��"ڝCËP��t옞�.~l �	c�*&[��c�(O�S)7�p�%��ex��dL�e��	��I�iO�R_J�/�^�}a�i��D;�scc��RL*����t�f��hP�t����2��9VZf<f��t�Z��V,Ckf�|{����d����&��%q�!��J�V���\f�P������d�$6	P��~\�N04
 �ө8X�X\s�" ��3w��S��.�tG≠��㉌m�!�F��k
ʉ(E��ł����<޹�	8Q��+����b��
�/�g�wN��z�>�{���_�����?�-�Z��>�9�y-�T�dЎ�زg7��1<�k��E |,��
X��Y�1�P���Ru3v
���E* IЛ���NE.�����+7�MM76�1+8"v�1"u�U���*lX��*O�pK�N��v)�V�0~Mr�V<*�O:��@2�?Sp�Ъ*�9�FC�0(,N 1� !����x�A:N����! 0P1��%�<����Zv�po���9u���֚�c�q�0լ�֮���e״�F��@H:���@����&���v]�ܼ��d���&PX*�*1�l��Q);-�V�V�M�:���P�~��E]�)&�sjF:�D�n�|����}cFL%���}{qd�:/�劜��X��.��*J�V,_�fu��šu^;�~�
����f�.�?m�_��?�ҕ����1��-Z�;����E������tpMI#�+�ϛc'�x�.Y�����t�����q�)������O�2��|�B���B&+�!�X,j�E@���d��������2����X�9M!��]t�m�.[(
tJ���99��('+}-�:	�Ӻ��A$A�' ���]I���E���T����P'��:��M@H\F��f�h�U4:Rh�u�7b�Me����ԁ��K�܈�"b�iKv���S������i�#*�09[�ߣ]o�<t���'�=:2��6nĮǶ`�C��F��L֤�S�DQ8C<%�b�b�E���A�+���+�%��y��
�&	�F�e�A�&G��YH;9t	�9�]��<yf�D��7_�|�1�ڔ�
��.�]�V&d�))���^C`�J[2X)c���Y;�ne�6�u�x>rQ���o�9��Q�~�߽My��@�<�Xos�gW�'�=�0�Π�d�[.��čw>��w� 2S�v��x�I���|� �9���e�����h��$[��=��a���,���|H+`��T�Do�@�!��y��ޘk͎������&�+���r����N�R���ܮb��d�az������߀=�:�궣S�d��@�;�u�"q%�n���v����0w	�:]�]y5��PŘ�n�Uhĩ҂$���L�7�R��U�����6��ϰ�
���H�j���79� �#�]�qS�������LКup+֯C*��d�&+_�7��L�e��m&��A�(�M�042��x�D�`�y0,�X�����)�v-��܎}۷!l6�uQ0^,�'8�~�o"�Ϡɩ�1,PiZ�|�r��|6#�gҫ(�/��y�YG��':���ZssH���s��U��d,.�K��@Bcv�bA�'�q����0͉)B�4F/��q��J�(1?E�ƺو�]7���)8)#��@9&\|�<j;��df`�2�����ɠ]����p� ��kiB�jD O}@L�S�!��@R�����\R��P��U, [,)�=�+`��4�X���x�Iԡ�;�J����g���/��](ضmd���`֮��p����Q)�1=u+7�ǳ��L\���D}f�B^����Ì����# R��n���:��s!�L�E�Q�q6��q��C�P�����l�l����Nk��L�r	�25E��il�Se#�@6I0×� $v��u+���)��נ1]Ȉf�%�Lu&��Xx�CE-�l�M� 	�@N�L�;��x����H_֭]���ᇑM;8����=Yԑ�6�iT��g�r@�g�Ƚw�m^� �m>��}��^���5O1�Z�";Wq����Ȯq4�Y��B�e��=��؆3��5�`��L1<��mOgL~C����[NOd�G���)��Y=?/�-��t41�/5,�I���q������n6�(c��E@2��[({-�0@�ILL�J��.�    IDAT����4-S8�m��I_���ؖ؎�H1�a�C@GǤ����Q����f��˜�8lM��`�yPlN�U���#���O(�1�|	r�"&&���&5��tP�����Չ`3c�j=��!8��P�1�A*��`9dqV.˥gx�r8�f�u��c�$ey'ͼ&g't;��Y)߭T�G�X�v�.
Y���ދ�&�C�5+W 擄�-�OA��������wn7`9)�Y���)���iq|�`D���#�O�T�J	��FipX���~���	�JC�dle�C�;Z��YX���Pr�r�w�y��<�i���ڰ-�GF�
|Q��mZ42,�3>6f�m�T�fј��v�bG,��P�WɅ�Ǘ427??�����}l[����,Rism�zfʘsE�!/'��=,'Yڈ1�0�F��uba4�BL}�Edyь,R�Zm8��#��ٓD���dS����ݧx�y�٬rs$�vq��'��[��h�Q��P�N���N�E]���03;��\��gb��1Q�8�)���$V�Ϧѷhs�*��p��رym�[�e�nxo˺9�D�V*��#T�)}F��٩q)7׶tT�7ivd�w��m��m�Xx>2��M���x�D����|}�{2�ڰ�������~A��	=p�Q��Ң|��4T)c��5}[}�L'm\�׼�y�υH{s���uv�������Bo���ީ�[�+���]qZ��z'D�ca�T?�w����9���ol^>��&9�l��a+z�I�-�L��|��NkX���졐K��sa��k����i�
�0��I�䐷� Ͷ�v"L�m+�}��ϼ�X���qm��BS�ʸ��flBI��
8��zc!w"�dG�����eK;���Q�U �)��0b7a�8���@8jaP�)Xh��'͈z��L5Ң���_�@�jhh�U6��f�-��lv��;H��c�ʕp�9��dW+MM�W�@��BwvN�¹��I�����b��]d�+M���p:d+X}���; ��a��P��b���L	.�pf��|�\����;��h7����N� �x��P$+a='u���*q������@��!�8y�֐�(Nn��U/stܺ��K�Ϣ�ǜ�����0)�>��e�99��!�]�x����S7��%�磌<O[���]G��W�\�'�ed��.�����]�]q��ab�NXnV��6�|d�h��h\�DSa�9:�G�e�h���9��J��a���ɜ����4����n!��ŋ�+��q�"��ƌ���0��I�,���)�n춧��kq=D�\���0�id)����s���I#N�<g�|*2Q?��;HQ'�{HgX�3��-J��q��UKQ�N�r`�F�ÓD:H��:J���!V.Z��]{ph�X���Α+�qz�(��t4(������?�/��;ֵ����{���8O��9Պ�!0�D�uXt��:��f�lQ��z�a�<>��!n!��T�\����j4+<��Y b�P���(�`EԈ��v�
5>v�ء{���xë^�cFr��3���y�ٽ�WA�V�\����.\��~;W`�=���4Z~�f'��4�Ny��'[���14� ���$�,�`wY��p5t�ߦ��	�%e�]ZRy<�tIB�E��\�`p��J�E>M�,v���c:�|��U�D��hz��꘩���[><�GƁi�1.��ھ��*ʐ����P�.R��d痤"n')_
������M�v�q^���~F!������旺���M>��)���N59��JF��0ޢsP����HC���}m$���9a"���(-����u�g1�r%r��]u����њ���/�#a���pǦ�;*�]����e8h˝��0%jg�^,��y����O:�
]�m���/�j5���)��b�(@r��!x^]у �B@�9Z&e�/_�y眍[��]L���.�S��Ug�q�
�?橸���L\B,ҥ��vv��� j]|8�G�uR��R�M9X>:�]�?������xq
œT�o�M&���
�B��5��������-��m�]K��К�������7�U�,��H�#N(Cśw�K��ʔ8�	�����w�v�!��Uz,j4	L���пhT��Z�����������^�W��~Wff}�)��׉��P����"G)�{�%8m�QJ�& 1���O<鰃{n�."e����G��3@�W�'"7��k��
o��M��V�E�����s&&g���E�L��q`�&Mԙ�����\�8M+��3 M5 ��W���P�dǍs���q�)���'�x<�8�i]Nk9=$^��x<�5�31_���&�
�x�l�z�G���D&��Ï<��܌B~v*#g���+�fǶ'Ю����/8�5��F<��z5�og)�۫_�
�.�_�"�>⩳ ӓhu���2�h��m��[�����VC�!Q��c�8��Mw�ΐ�LQn���5�r�F%��P_y7��#�ڭ*R���!�[p�"�O�������Z6����50Y�`r���j~"������A�9$��x� 
���fzÂ��Uܱ�L�����t�� $>���%E�(%d�PZ��� �B����H"B��$.B$��v
Ai:��s��I��H��]��H�0����;�Q����Е��B���l�*L���I����i�t��B��wuw�]nǼ���4q&swR�ҥ#R���������c0]m����LH���b;V3���3�P>B��E��!�(>�&�rVT�N]���/Q���a�����9�sv?��LV
9ieT|���#ݩ#A���&q��S�}�����F�`�i��"�R�m��h{8�������135o7� NiԹ�L�O4���bI�!h�$��x�Je����G�R6��_sLq�c��d��y��9�,�9�������x��tLStH�)9���J�d'�h�tMp��
�I#�_AyhP��Z��tH��y�Q2m�S�kn5$"���`3"e�/���FBI��wI69�����m�����+�����NA!e��œ�l^;]�Cxx>9�����D�K��z�s��(�h�37uL�<�Y�aρ������hOO�#� ������pxsȎ�O�X�p�ݪ�s*8&1k�)� AQ�ǳ�;���7�p�~�� #��`����d��6N����d+�Zr���������4P/�����}	��n�)>��C�*"
������أ� Ex�E��SWci���`-���g�j���㽷��a+лx~�Hos~�+�k���Бq�IGb�2[�α���Al�ysA�3��*�n!���G'%C�;�/ii	�+Y4���4�s|,��d(���a}�,l��+���41�_��nJ�̇g�����<�}C��Kh)�jb�E1���&0Um�'r
@�Ug7���1���0Q�P��H9u��\VŴ�%,2��03���ml��7�6.������ُ&��ߨ�;��-ь��%̗ᓱ�):;�f{�P���r��"�僘��;�<6�5�T |��j\(�t�jT[4}��Q,���И���;l�M�c�!,�E�ˑ�v�:ג�TJ����ox^*Y��r��\�a�kq3 ����wy6�����l���U�e�j�-w7�C���|B�)$�s���	���6n�e��,�ޫ{uu{۾;[f���7{%R? 6�=G�Jڽ�3���y��}����d8�G��uqo�m)����d�G�����K�y��M8|�C�D��YA)��Ģڢ�P���t��^:��.\�<>,��:���,�I�����E����7]�����۷cr�
�cТ�Ur�raS���a1���4�j�D�M8̦��W��-��R�J�����	�O'Ë�U=\?=]�D�K^/x�)�p��0<�$����uç�\����"C��ՄR�t*���)�T8��=;7҅H��y��P]B0)Lw$S&
B��g�q����P�K��X�|�Z{���1�IW�N[b��')� �x���xg��ۑ�Ia`�n/��E��[.ڊg�}Vl��ӳp��i�PV�G�Ϩ�`Q�R�T��5���$��R%-ҼB���\�H���!�Oj�tCC�0;�������6����H��/~�qϽ�$�T�Q����]QQ�2T��'� 4kzg�Sg��&��������
9u��O���02�BkG�L�V�^# q��cH�Cx�����5]�I�lT
���5���-�����h\<�����_�
�3�y�ʶ���`bx:�{;�C�I "B�0E�ٴu�K'[	ym��W_G	���>�-&�.#���t�����t�� �K@�e�P�g��V�H�oԶ]�����\
��i̤
h�]��f!�)atz3E,��]������~��g+���
C޹�!i�Ԅ�A!:lv�Y@Q#B��4'U���=�����b�wH���bs�Q�TH��	H=�0DY{�I�'�X3T�!�`+������ᒫ�A�88�q��������+���������8ji�2�S�j}zD�O{۪�gm��P�̼r�҃)���v�[Z�1MkX���&��z�y�@���V�t�4mO�'�mI}W@Q�&T�2�)�L$ '��ҥKP��O�DcDm�~e�H�:�ER���@�e� +P%h�3�Q,��z��-kV#mg��$�f*�5W\��ys*{D
?���X�Z�3H���V�=�%�4'�
W-���^h�"��x���Ә��\�ڍG�Qϩ�W����C�3��< ���[�G�VS�X8�U1nP_ ިP.���6��S0]"���`V�ln���IA�S,8v�%�[]/4j77�_�V@� �v�����
QtE����+o�G�F�4aEc2��"��\:��ڍ"��0�z���p�Ĉh{��9�˧��ω5�aX���)H@St=9כ�`���XѾ$�G5"� �@��!R.���:�R|��^�	�=�w����f������L��4��'�ܸ��C�g�D�M�j�D8��e����\y�_�3s�(�|�C���qD�:ĄdŊUB�D,`���.ĶW��%����Z¶+.k�P���p����@���_r����[��C�lj9����ޡ����Y@�f�L�����x���,�����y�Q��]MX�ތ6���+��aE��C�>5fYط�BV�!Y��}.J�=�,W�~�p��Kп|��s.`�P,V��O~Y�K@0с���B���TSsE+�]���h=��*�2�
S�J�� DҝY�$���V�pCQ���_R���?'B�2�X|��Sc���uz�wO�bL��UR�(��;-{8}�g7^�A *��J�fw�*�zKf".���-' ,ٵ�39T�9������x�{J�p�8�K7a��2�h��i
��֭���T:��Vv�Y�8*q�ș�Э��2VP�j)&g����-��FM��N>R����M=�~ug�E���
����eA�Մ���ގX8����1q���L�YsNz ��t� `Z���[h�������T���TQb2<il��
M�<s��������Չ�5:|},� $d*�6����W"73���������Ii$s�C��I\]`^_?�l�u��4�y���&��u#���I���N$�N� #���59N���zw:��U����L�l����ҝ��S�Ms
��Q��>�2!v� <��h5e��:0� �?�F^ ����r_%�{&���<E>�@-��2�O�F�f�j�������qrĭ��o�-	ь��t��M1+���@jm����E����ע�	�sQ@�wr{յ4uD�.�rz�;p�e�QH%��(͉�n�kǲ�K�Z6[�e�*����U����A��*��I��(<����y$��ak:n���c��G��0��oI�d�=�Z�����x���cӊ��i�\�U/h$���W5V�_�@�4Ί�
���'dR(�`�\�``d����ށi�U�)�#=�)Ĭ�	c� r��a��$.\ߋ�fKc!�_Ҋ��ތ��#8������m�\�Zf�T4$�NUi8�ժdv0W��İ|�98����w⡇Ã�>���$"mK��5�m?NNd��kH�*pHYp�mw�SNJ�j)*p�ga��2�G�1J�y�էN�s���ǯ^��.j6~�R�X����W������C(��d���/U���Jy��l�E�^�{sZ!	�^>H=��E�T��ز���� ��#�L"hXn�9�m��Fk�h�|VQ8@'ݨ�Q���ՅZɑ�)l�Ҏ�u�
��)��VP�/s"#����eǛ:�����*��OC�40�s3�b���W�E�.��%S&2�R"E-`F RU.R<7yM��������ĸ�ً �F�ۓL<�C�0�[�6�9�ѹtjF �|VD��X��	I�O�`@�NI�� �����I�{f�G��:��"ؒ@�(��jk�/���)��P`ҧ�~Z����G��R~N�N�^�g� ���j��Q���'U�Zk�<ڒ���У� ��`����u��3Qѯ�vE A�[��
)]�^�W���X����6�"�����ݸ�i�p$Pi&*���,~71Ń ��UO	�tS|-�����Ѱ4MH��Y'U���B
n����,A6�K䠀D[�Ŵ tj�%�ׁx5�>�mFq6 ��*���1�Lj�Ji|�����.E���j����)$��h�P���yì�T�zOjX=#��&i�.V�%���)��p2S@(ф���W��}��w+�*�tk[�L�&O�B�q�6�����{[PMϢf�pݵW7j�F�X���
4.����5~�7w�ܳǭ�5dKe�� ����BYG��qI�"4��jѨ�Bnz����;���ڂ���f�훟x���X�o�Q���
U\q)�r�hRX^�H���XZ�R����	�uox#K��+�O~�f�p�fdmR�B��88qr�D�BѲ�@�B�B�J>�	�L��r�UbZ0<Ͳd"���\��V�U�ʭ�畴?'B�$�L;^�&�`�Hr*�\ �uQ���h����X����8<
�t�i[!��Q:A1��
�;W�D2��5d�������G�t.�v����S�~]!+���`�q˻�%<��n�>���
$�[[��$3�Rq����b�V� )6�ɗ�OvT�]qzN���W�o��������Pⱡ]nݶ���ynB��xU�X�lN�8!�dYA��`СA=J&Ƕm�kePd��x�E��*z�;�M �@���P��2�$������htHz�Or�ڜ����^�,^�{�x-��9�p[+
^���彽X�����Uʢ�8�I����|�R�ģ��"��}5`Zy�8��{^�J�b]e�P�N�ʔ��YԒ����3U�*�P���ޤ� �ni	)���.6ؤ�쪄3���	"�����ɐ��%�� ��E*p�rxy2��B����{��r��ָ?��J K�`1흓4�2�>��UV�p�Ӑ�
�T���q����Vn�n�1���H�DB�;�Ś�@�����S�]9"����AD#-Ȧ�Ы6��*��ُ�%$L b)�w�T-	ŕǝ����60�uy���H���E����u�5Y�_�{�fR�k�v4��/w��;�k������B1_���(h��m���߉�X ��|�b����=�5�@����ϯxf�~��c�.�X����4�;��'���,��Ƥ�9o���+5X��ji��ƒ�Vt��˖��붢3d�����С� �P�Ё���t6#�����fʼ��Y,Z+*#�S���\��� �ũ��k֭G��s��#x˻�#�	[#W5Qv�820�\IC���N�֯    IDAT�(7-2�$dСX�&z%J��5��
�Z��:�� �����,4�(S�@׏��	�r��b��+,:`�' L��KkbHZ5E�5	�[�.�Dq�i&Ģ�K=��ChD,J�t�
?�m&��6I!�"D������ ����Sd.��U���]��9���q��7ࢋ.��?�{�K�AK(�l�����)xeaƔm/{ ��K���u#�bY2A�g�ӈ@0�c������'PL2��E��/Yp�νr��'@L�T�Z�1>vJ9gUH�х�U�)�0�?d]��ʽ�V�J�$S-�Vn~?��f��[�-�me��Ae�R5Z�J�&G�j�r&q1&�&^����	��^H1K�@�ZKѶ6��*����biw7���Vt�"��d�|	�<y"wqR����/����DS� :��$~� J ��ޭQB��v����  &h�E�^��Z��zRIܴ�����19�Si� � ��\d�ㅂz�9�A��y�h
q�EN-~݅�/�c���v�k��#�p<�h�%��@�l^\�L+���m9����� �25Sb{i*HH�0����8|]� �һ����Z(�Ke��C8�����#������e���4p�]w�%�TIWݐ���Ⱥ.�Wx�q���s�̠E�����1S�<>�s��48>�O��x��	���[&���P��056&�����?}����aV(f���m�Pϯ�{ck�C+иx�C��)ύxb�n���ݔQ�9z
�>��C��#�b�'�h���B�����SXݗ�9�q���=o�MO>pv�|K�Z�g���cN�l�ZkW�e�͘.J�p�|A��`����V�B�7r��%���ۇ��n\�p���Ο>
'�@ ܆ٌ��y��2r5�t�����b6=�_��D�zg�E�a�+x��S�{�$D��_^(B�H[�ԟ9��nHgP��u)8)�e�y�NT�N8*��u���|N��/�j
w-I�"���A�#!D	�bQ�%SB)	�tq�*��[(A�t8����;̝� �#N'"����^���]��۷�> ��Q��xY�!V\�H{�<��n2�*�����`��«'�!�Nt+��p0��)!L^=_㸰������+:��߳J�.�,���9��\0N�H�'�J�3~Yf{�E謨,%N��w�zG�]57#��&���a�T9A
@���O.�M4�롔�M� �]fe绘R��MdB��O���$:ڑ' ���԰z�rL���� ����"�_HLz�wЕZ[Mt&S�9��P��H:�
�,����=�S����՘G'��ɼ���#|x�2��SO�����%�OB&��͢�}D�Ew�	��H�)���օT3�1o�'���W	pTz(�C��Pߣ*rX�SsB���mQ�T�h��=�(�N������ɆD�vQ���,�*�!AZ��±���*�7���P����-�yU/4Ne�-�Dt=�i6H�N8������I���o�+o�� fgS89>��9�[�(��4����\�q����R�'{�t%�V�:"�!��b?���x�嗡�%$���������]G������݉b6���1��V���ͯ��f-� ����/��QC=7nۍ�x�@��y��&��V`p�;F�<i������,�|v
O=;�Tɀ�2���	�P�kh�U,m����(��r.�Ѕ]s'�ʎ��v�2�BѩTH_0Qrj��F�I�U��(�N�Ɛ2ĢY�S�PC<�E�*�/4�H$�J����b>Sě��.�m}��W�����X'|�f̦L�JHfk��cQ�_W��R�r�@j
���H".s�����"(Ű#�/��R�x���b�(-ҳT^�@��/#O����*@�6��K13��Y@��TЃ�e���F;S�p?���:ۅӞ�md��ui� ���"�g��T�l��.�۬a��?~������Q�wbiZ�?dI��M�g�DHM#8%I�W�O���h8ҥV�<<{cfVk�
V���5�194De�z?Iq&��l�v=M�P���$��S�������DxIz	�_�B��7{��( ꏄ���)�0�I%*��R��0/��h�b��p�N�<�<�'^rܼ��b��Z�P�ҕ6b�� \"��dkÚ5��ر�2U
E���sOhU��(j�Z۳�T��e����#�ѡʛ��<V�_�ר�d�^9�)�I`�5(�vZ�2ȵ ���[��)�T�/���V��>�Qv����-[�ݿ��z�g��y�����&z��ʾZ	΅:XVT3:�	=�Ǔk,�^��ͪ��s\?B��OQ՘�N�N��3ļ�:&R0�= �|	!d�B�L0�>F��F8*���z����&5�������Z����mn1�W����Z���/��@
������G���a��l;'z2գ���9�t�&�1�(��~�.�tan[6���n�
�<��Nܷ�	�g+�P�����F�����8ly��Ia5=ñ�w��_ݭ����V�@���.��V��]�\:դ6�EC39<qt
OE��K�H�!$��)f�ѓа�#�.9����Zu~���O}=�1XzPD��wO/���s)�a	<��e,�@sK;L#f7��a�(��H.Labt�VE<D,D0���%FR�E�8���q�K_׊�K����h�]�|��l���0�v���f��Q;�|RPS��0<�Gtq}��T^��`&�G�a�ر�+Rn�L��Uǔ@�)�yF�5I�;����ְl��D։�|of�hb�	k8?
�u��É�t���пy̦�f�$@Ow}i&�$j��ʪ�ue�Y�X��A�i�6��~̧>y��D_/Rɤ�����KR�O6T~�q�4�>pHQ�k�9��u��AVw7
��>���uu��(LL����t�a>� 
���pT�U����"(�mu�v�ɓ'=��EJ+�
v���5Nm$������m�R��s�"	�b��Cnf(���9�דz#�L\K5U#h$�_�>�8}��Y��p�hg	"��-�;,���}ntcG����W�*�A�JU�i�LG�:���Q�ZY�
U����2�P �y=u�(�Q4P#�D�Ջ)kJ�(������]X�+
_MhY,�	�$���u��N0�4[ȡ���m؄�ӷ D@���C��t�uv�^w�zsI��h�2t�N�T`g����|?��9YU���Sᢚʜ�k�;.���U��f�A�(�U!����ټ���;��DE���K�m�˻��X�&D�Q@D����Udt+(y��V�X�7��x������]����G�2���杪�����c[���'��м�e�LK�	i�[.d𞷽��,~t�O0���5ð"0�
�ع<�O�B8��U�^����U@a�j\ue#��vwm����W�@gCc~nH�bg-�+"� �Yl?8�}'f���Qb\s�FL{v`�*3�pu;�ۼ7_�+�,?��<�!��dA����&3��t�J54�,ê����ލ��n�-+��5��=�.�L����qjd�\�RAB� ��hNE@L.WF��5��7czj����dE'���t���BM�h�����Waw RkX��
��!�Y�c�Z�K�-�Eb�j*�v^ɭ�ȭ�B3�ʣ��]��RZ�E$��tq�8ot��~ԪH1���^�#���2lP�H�	���˖��W017���5?�Rv*%t	���|�Kx��� �t����H��0B
ȩ�)����N=��U*Q�wEU)*z��@�s<b��P��RV$$bt=F���/����V���Þ��DzrA:B���i�� $�̜)�	�To�(�7��]��������O?�L�t�C�2F��L4�����b��_P��qar�P*�HA>�;2��AC��0�$�EQ��ؙ2��B請��9o�V�ӁLt�b]��2N�jx d~lB �F�9N<�(�2D$���2U��iZh)S N�<�����"0��e{+^�t�b�x]�����sJP�)ԧ�J��T{�& J�̀>�ѯ�a��Xg��'��
��QlZu.��97yM��n�U��SV��I�~�f�x���W%mhe������8L�&*eZ�+�*��t��x���P�S��AN*5A�ዦ�ޜ�rDj_B �}�L�:;�%P�U�/�d�[�d֧c��(}�?2E��ze� ǀ�� �����RB9�Eg/�&�E���s�� ٬|�;<Ӕ� g���<�yR@�&`�@z��^TJy�@(���߉t73,�_;���Ĥ|���o���mD`�@�@�Cc�V�@��񫿙+�	�t���nap:���8���s�VH]
H��.�ՠ^��L�M7]�w��*����n��{詇�d����0�ΣP*C7#��X�i:������4ݑ��݁��ph�^h�<"�2"�&S��m#������݃Knx)��Ç?�Y��nT|	�ϖ0����h�+^���Nn+;� eh�yev�����ÂF8=��>R�:=S��3D{�P���A�Tw���kB��ۖ�� I#%�Ž�����޳,�5������bh�|� L�40�z.��^Ȉ������(.,�XQtZ��%�E�P9j0;Z�[	�110$�V�p�-J͈��Jf����#�^��O #��ԐH��}����;�%��Q��h�%pުU����=6�p"�|*�-'2UtIc'����>L3(�L�6CAѽp{B��d�Q��H\�T8�:�t�2$�Q3(�\�/,HƢ��ɣ��K=sR���K���?`z�r����] g}M�i�k\+q\�]q$�H{�2�p�j8o�jLc�� Gjj�%ZEKb)�}���W	�|:�Sj2Q*ڲ�&m�]Wև?��Jp�Q�<ᷢ�p���2�
/�n� �q�ǚ�$jTh��cb��
�7�-4�$$C�nP���ظ�<�w�OdʢW���D�Bq�����O���p����D�@C!b5��Q �.�7�"!�Ɓ2�౭��DG�O�2�*�gl&�[Y+��@(��%KD�N�Z��Gũ)w�r=�U��˴��c8\;��]b�L���I��xCEM�)���ۃ5k����$FFO
0��J֛�\~y�	�����z��V(n�8j�erO�dS�uD7V)ST�ݲ���#���i��t$,����CS���S��-��+�i�P��e@c�~+иx~������
�=��"/�+�����:���=x��r������j	F-��@��Í[��vo���{��X�݊_�L�A�\C���7]�e��o^�<�}w��!$'�����Jh��a!��Ud��۲kο7��w�޷������B-�����
�XP� >>\�;>Ts�A���X����E�*��a�4`��R�R<k�^Z	�kL~.1��D8��E���@��x<�J1����
��sRh��A���ca�ż�-�A.�@k'����o�0:97��-v�&5��4�L�.�
��7���l�� ��"�e?Z�F��Ƭ��pS��[#ԬJ���#G����)��ϱ���fB���:���X`�\э�.6J���5E#���˒r�@[���ۀ����1X�(*�jN�HD
1�=
�>%ȱB!�1���`8(���h>v�k��D�Y$�r���hH5=K�ѿb	N��"Wb��)�|
p��I�����
��d3ќ�h$G�@��O8-�V ��'�RQ����Ⲭ�R(<nmAQ45>�֮ũc�' �Ƈm a��Ge�¤,2�|��4p�D�2�(�R��O1g��r�*̿�i��C�nY,�%#GM��p�(����7UN,�2LѺ�Q.Zf���l.'�4AH�S�������[�L'�v�ɞy�gO�������&�+²�%Pb�J&5/�t�X�m�YIs��DtJ��tb�ݒ{�	���8�TF��n�S4��� 8�Q�.�Ӹ�ϳϕə�@�L���D��IA����iw[��&�y)>?�Ѩ�@q]q�cs�@�%2R�=ұ�ϑ�o���g�Q��hZ�p��f�"�g�T��Lg�3����d�,0%�S�qܟ�_G�.��Nsb�k����юJ����	����� >��7�ɪ@�S0�
���?�<z��[�X�_�
4 ȯg���<Y�����)DcaрT�A$�~�� v���B�/��9�N�@�mH��O|X�q�?�{�ߍ�x �R^�#E*�"S�p��߂��)�]99�z�~t&;���c���Wt*H�e,?wFg����އ����}qLg}<�C�b�XUv��S@��q�Y�10�� ����k6�c�G����`�8�bqd��M��O��wa�dS)��֖6�v��'����n<�-,�YS����i�����p��/C��n�!K��Tr�LF٫&ʚ�}��H*��|H4w �/#�����b+������W݄믺v.�o���ؿ f�IOIYq�6�*ԟ��N��sV"��])�����āC��Sj��;����@Dq��u�'�o�{��vKE��E����n,]{.��
¦�-7�;����"	Kǟ �p�Өs9O��9= ����n�6�T�,9�Ш٨�e�â0�+@g�\������.t�v�X-�������oݎ��^F`,��8W�M2�P&iBeh��`�a��J�DA�2J�}��|aeB�ĩA4�`K3lqmR�\�_��#�0>pB��eZ(ӱ��RNr=�:Fkk+V�X���� @3�x�6uW��O 4T�!�D�!������,6Ag0+,4(ɡ�CUM�j�3�,�RᨿZ�l	"a��ةhr~W�N��cT ]�X��������m0[qWF�rvwo���"���СC(ХM�҃X�|�t��H�hG!CP@k�
��eTs%�z$���� M��Ϗ�X��槧062����z&Y
z�_"����s:�Y�H%@ Es[+B��҅E1��/8� �گPHhs��QKC{j�v):'��nVa���}-��ue5�~VMC�R��#A�oqj�s�����T/�F�{��#VT=�j:D��e�}�g����u'�޷��1�RF��.�z�/��yr{llfc~�+иx~���x���
<��^����x�b	)��|%������y��٨! 2���&�їp��˺��W_����ETfF����b%��dtt���U�|�/��;��n��)������" ��쩙���L@���`6O�j��/cr�+�T�i��m	.۩����O�6#lq��q���܆ �JⓊ�CUg����St��W��2\{�՘��ſ��N�޳��6���	r�R���I�U+�7����+������3�&p���q�C;$�=mA�� �S�?��,y�.�`�%����p�����X1�*� ��i%_ ��t.]�t��<��� �u+W���H��-g~��5C��X��PE8lI��S+�B�0(�W�<ԃ�r��Ɨ��-[��ڄ��Awgw�p;��#��Z,!�H`l|T���NeY���<f�H`��5�l�D�@=��0���]���k�-� ZE�Sit@A=Djv�~ի�ݯ�*�s�v�喦=66�~������=���z��X!����I[	�gL�V\!RX�N~r��S	����fDQ�J mscqX-q��Vsp�ƍ:|SC#@ر/�	(H����)���8ڇ��\~��ػw/��=+�}�p��O�X�@�\D&�B$B<��ԔL�6mڄ�	�w�H��K12|
�c�w����ǇN���*l��	\��r�\�O=�;�? ]��B���C{{'�{z`�6z����}K��qWu�˚��ȓ����169�T*%nx�t���˵���8�.#�h�	�����`�a�UG���Uː% �@NV�_u����dx�`Vz!��&!����[&t7��Y4��u��Q�[2e*T*��~��d�!���ԘB!�J�;�Rb�    IDAT���t���Кض)��BQJ�S!��B� ��}j����!��Oǲ败�Bu@��Q�v�k����1�I�C>S���)�U˖b~v�'��9X�ӄw��oaI�����j�<�o����]���f�?�u�o���y:�N���"UƩa.W�d��G���ɤ ��� ��E��E\�*�[^�	�� ��+;���.�t]�6È�c��m�_��uM���Gz�$�zn��B.�XŨ�l*�[>�|�o��{ݍH�
��A�M;�D�D ��<j��mN)�e�����7߀�����ܥi��������y��z@8�$#Т.�
�fp�K��{��f\��C�c��3��p��p5KM �_C~nZ��O}�V|�m7�kgf]MWV��&-o�^��ɖ\�o`YP�vNW�������!��H���Bf$�Rr
��܎��+��^�&w`x
%�w���I'��Pl|�i��E�d#Ϣ� $A�\��u�1�k/�G���J��|�34��֖�Zv1���iZ,�u�OEbaLN��-������D"��[�bYX��zb�����; �O�O�sJ nL(�%5�T$a=�D��òb����K�bt�(NF(���F�.���"�����ȟ���pw<�(�{O�|�'��9�o�@vnE<�5�--T
UD�;���%�NL�'r�U���5ѳ�S�e@#}�)�E�,�*�n܈�g�ab��Ǭ����5EQ�d4t$1�Z�J��ȳ�0;;-T�x,"�U���2��d�:�Tzm-�t8�`�L r�9�b|lM�&lذ	�n߁]��b���M��û����˶a��^ĭ �{ڱa�9�eS81x�[�2��v�"�G�f� ~����Q�MM��ȑ��B!\x�Vl޼Y������lttt`��v����U�X+��8�@:U@�D��o��A��?ꀊ6�R����q23>-׬8�yB�z� �����1��'��\�0��~#A���J��$�n��M$�	�Y���T�tD�R�DL��(�job���:_$��Q`O�,�vJ��Γ���&d_8��u#z���lbi-�tW�b�!�h<o]tt������9LPo�԰�����F��0*9�"�����}�k��5>����+�  ��������
���#�F%�
R�*&2?:�#�89�V�F�y6����K�6����m����ΜDsʹ�L����p������[r�09���HM�"5;?�yOq1��^�����|�s_�m�Qu"S	���9��Ԩè敫;�bXU��f�;��k΍�v��]�[߿z�G�!��1�ks�A�y�TZ��R��w���.^� �t�]�ah��׻�BVS�<��5������W���_��ω�CV����M����o߁��184*��䎳�r����3g��M���{�#OI�t! �j��x��~t��}m>�E�G�?)8q=�t˅���g��^�U�	A��==-����4�" ��_,@�s'E*����}Z���_��/���;wb��]��J��݅��1�y睘�֩)Q;;���H^����{߿[,eÑf,�- 2��k<�ླྀ��ݭ��4-��uK�K�ŗl����F����v?{��L�ܓ�t��1�:5.ԗ�W�T,��cρÒ�rl`P �kF�PEkG?��4_N�T�39�g$�{)���E���"01 4?��]�y3N>��C�ߒi[��;3�!5��+�w��w%��V��<,,,��]O����H��bddD�{�|V��#�*��ЃL]G.��d�����]v&&&d��Ҏ�� �΢�Rl�r��?�w�����tu���P)d��ׅ��&D#���[䜻��+�gv�!V��eۮ����qrtX�g�hK{����
���Wo;=s)�>p�>��O��Eu #�$v�S)�u�r����k��-nTut����x"��t��L,�@Q�PP��
��8� ؕ�ʊ��L>���[2H�"�&�;'"����V�h��������u�����\$�D(\�ԁS��%q��t�.8���?S��i1:�_����h�$�ݔ�Q�}����.tu� 97��1h�*V���=��
tD�N�W.��������k����4V๲���r$��Y�Ǟx�e��yW�LAÎC��H�T��ϣ�]�Ҹ�_܏��r���O���h�L�yX�&�h]���^3����E�����1df�1|tfF�����WE\��Zt������`h*���s���Ϊ�?ҭح�tS
UV�Z{v��:5m�д�q��f������$�PA+*�7`�𹘚�uW]�n�y����~���fͷ�J���ac�qQ��?|��5��cxf�]��z��)۝��E�PE:WD��˖�bjl� E�>�r6��9�?y��k��ѐi"j�{����L�]ў��|�}ƽ�����Y(<<�ys3:��a�BHQ|]�E�]���V���8�Z���8l��%�����~�	� U,������Q��#ȼAhom���R�$��zp�W>'���w�ÃC:��{w�ȱg�hnFs{~�U�Dk{;��(���#�=��y����\��%������W�eY��Q,���׍?��{�~xn����$�m~.���$ff�������֞���B�/��%x��'0rbX�T֮]+���nR ������|���;wx�&�W���iN}"(���&=���,K�!�n�0{J�NA��L�pg;�U��̗���7c��̍�
��+�ZL�o>��*.ٲ����	����	�:X><:�r�p��A�ڵK@���T
�jY�bs��afr\��׾���G�ؽ�iD��@^���)º�163�;����T�Tl���Д�
0��a銕��g�C�Ś`#شy6l� �ɳ�B���m���+��k�.h����}>�7�C�XBU"n�ό#�)é�p4eAK��9��f8����($�b�y�T����v�����6ԧ|��1b�	&*Nv����(� Պ�6�VĻ��٥@���P��0S�P�ӽ����yZ!Q��G��Ji<�y��޿I�����y�CV�����_���d%�wkԥ�h������d
�N�@�0���	o}�K��'�JjZ��믹�QC��G��dc��h\<����g����S����*�� r5�d����H#Y��h;"F����hu^rQ?^tA{��3,� ��4�@��/Ök�Wz����f-���Cx䞻��ʈ�x#��L
�Ƕ�_�c�3����F狈u��hšS6�%]��TPX@D���G@+����o��\mx:�~�xGg\�|+�}pj� �Mm(�T�E\u�|����:�&d����?�a�݀��M��f�
��%mx<�.�	/������#8�.�"뚞5�/U��z�����_}���0==�eKW��%���r�[�B���Y\�i-��g�Z�����?�q7��t�X
��::njBEsQ��aH9��ӏ$hWš꒍���g�#91��
���AU�JX�Q��-kq�U[��GS8��k�`e_�Y۱����'�D1[��l�@>�F�.���Ø��F0�%�^�o�Q�v=�$�F�p�׾��Xv���ǁ�ya�K�q��g�f�R�Xڅ֖8.��b��=�G۷k�����>�S��W�Y%�v��8��'�l�R	�;t� V�\�/~�gm����;߻���xv`X�ͭ}He��8�X	����y��u��|�+`�5����GBD,��������ĩ�� �Xt���{��0|t֭j����_x}s8��ӳ�>+ӑxs�-��h���M�C��k�u`�~,�����
2��H���FJ\ή E ���&����[�b	�� ��a�*5����{�Ǫ��q�ŗ���%��g
�`s3��y�V�> �Ϡ���_~9������_�;�_�
Ʀf�����E13���
~��>]�YN@(��l�i{���f�42��tQ�&�u
�M��bHkS� ����ūߕ�EϬ�1���H|xY.`<������l���-I�kE�l�@��V�z�� g�c)�{��&+y~<���^��"�������! ?'��/�����͹���+иx~��nc���+p��1wrfZ�k�`��& �ާ�
�X`�K9y\��/��K��:�qVv�h3�+.�/��_�u6?q��;9�ғx���"�[!(�i+KN���\���%�o���w����H�Q��,��I*�E7�Y&��Wo�����*�i'����θ������7��|��(�t��o8w�������ȴ{�R51y���{ۧ��G}�����;el\ލ�~� ��伻��E��y��ݙT:�t^5-X��(�+��E�����?�;^�Q;�-���$.Zڭm~�[���O �Ԏl2���8N<�ݳ������ů}E
Э�8�--�Yrve�e�+�`Fe��3��b��5���(��(�Pl�h�����۸p�\y�z��a��u��u�~������AL�M�uk,A$����É�&�=p ���pZP*�Φ��}?�������b6�F&[D��
�D������n��|G{V�sZ��1<:��$F&&��݋��.���e���DH?5�/����w��}�ؗ>����'v�Ht!���cْ�@�(�TU�Z�J�(֫b���R���a��6Qu��s8w��>?����q���KP�g��?��\�_��_���=<8�>��n�SL�Ob>� �sL$bQ��v5z;���.%����F�c~rqӀc硑�
��X hJ
z�q�RGt�)�BZ����܌d�D-�Ib�kp���v4L�. BJ��bavǎbbt\�pSs�(q*����nQ4.>���/���2�,�M]��mH�\�۸5����H��\������oz IMG$2G]<�+_��x� �0��)��8��Fy�5�����B������z;]Q���.vT�& �(�Ɇ�JX����rT�gg���3��N'��[71�����/�~��,������ LM�ʞf��旣3�G���S����5& ��l�+����0j�rc�o+�o�aw6� �H�T��\�<y����r@
�0r�tM+^|a��S�xQ:URD�1q���ŪͿZ����#�[�EԬ��ށ��$�@M� , (R��]��\���B��|ч������N&�(VX��J�"B�.äT}���^�ݩ>����'�r;���V�o����{_.�)�&�s���g&3��߿_�Ν�b����Zn�� ��_�돟�rW�ujOM9��/y-B�}�����"k�!�afa�+.�U��މkV�����5����v9�sG�=�;�֯����O~ADҾhL
�*�j.J�jI�P��u><Y�r�V����wáU*iCՊ$1K#V�#�di����cù=����m��r��}�مy��s @8h⢭���I�2tm�5%���O�6��a���у�Q�,�W.	孹��J���.Q-x���J�,���҆t�F�T��s�F�6�/����'�M�e244$"d^L͎Ģضm֬[é��z~�_u��û��ӻ��#���B	,��h�4OxN�+z�-�P��6���`�	�L�.�D#q�4���;��'��dSH�Lt%L���m�ȇ���cC�.�����"F_�|��:���������X�z����n�������{1}r�m��5T�Yъ�C!���&i���0O�42;����L6���>g>[�u7ތ+nx�v��~��5����W������;16�(`f/�3B'�孷`Yo�����;��_�
F&���)�l�,nnu "��@ ���2Y`X!]�8�"ȣ�Z�
�Fx9,� ��z���� 8A�X���)�^������%Ĵ�nv��N�Z�`�@$D�=��t �\{g<d�@��'��A<��:�g���jL��N]��p�h�L����i0��xi_�\�'N �jX�����f��j��$��nxaC�|��7���� ��9�-y���#�ݹT�a���L'f����8xr�e�J��2.]ӌ�t�ט���0(rdȗaA�v����=��m��^g��\T��l��|3c'`.t5�xf���[пj�V��V%|w�Q/ ekRܘFXR�M��+����p�Ļ��J��i�ށIw�.���~�K�D�`c�n��e/��/� �t:����k��!~��cH�L4w�H�tk����0��7���)wU��2��h�n��׾�D�2���GSse�@�*" 5M�Z��}�j�F,����u�ԍ?���!޷Bh�L]�!��}�Yk���|����>%v�z4&��<Ύ��琷.ŉWI�Ĥ檃�7m±=�01!���JY	�]W '�g�� [�/�[~�X��4@:����N�.�p�� �FO�9Ź笖L��7mY�恡AwՊ�jJt�����
j�K|8%��ig���F���(�B.%C��5� fSY�ٸ׾�e�	��*,/�͋�/��?�)�ɤЎ����[�a=V���˖`뺍�=����w|�O�k�A�&�]�M���r/ N8�L-W�tv��H��j��x����	J�Mq�ZB�)��]FK[;�;�᫹xz�v �F[+Z�~��+���_x}��rG�O������Q���ߋx<��%��t$��
 �ʊ >�p����	�%$���JI�~�����Ć�i�TN���ch��rpA�*^��W��_�x�g.�7�������6i'Osw<�8��=(NO<&�g�T]�ᵯ��7*m�?~�;���:r�H+B�$9i"��@�L�(j@Bu��f!M�33�@_��p%'�����[� �:b`��r��{H����/��<$�$���PC�o�T�����yQA�̳��L��� f��� �L���6�sA�v���(e�LI�o�G�|I?�I�����u���7�$ �V�C5��K�k ���m��	����F��5il���8:8����B��Q�c6W�X����|{'�.���
�����5q���R�P�Do���+ށH��_�u6}�[)Ρ#a�ɝb�� �n	v+�%	���.
e��G	ʰ�7;�oF�ώ�b���5c��Q��2��*��铃X�������}/ݢ��sC!�B��l/��^~Ӌp�E�N/+��x
�~�Hf˰������\jKTR�ǰ���!������ڃ����>�u����tޖD�R�xZh[u`�J(�|��J.��&��+H�t�#35��/و�?�kmxj�]֩�]���q�O��3Уq��a�(n�y���3�M��&]i��ɥ<ps�&`����ԁ�4Bbk[��\�m~�5/Ê^��p��ĩI�؉Yہ�A��It��!�Ɨ���9rȍ�#��Q�b?����SG᫔d"f8���ޛ��U���߳�}�}I&3Y!$!��"�AT����.��Kժ�Z뫭��ߪu�*5��,	1!$dO&�d���˹g?��yν�	��k[,�����]���߹��>�w����P��(0Hg�h�C�Qa�,�_x�����Ա}�X��TK/	hbG�i"�}�v�#�?�}[G���Xs&N_�g.[.|���~�Ol��Ӑn[�Qm�m�=��S���j@*�Qg^�*��9ty�s��Akh�j�d.�XS(R�;�b�j	�����d�7�>��<�����g�B��b��!e�$I�����kYwC t���F4+�y��}O�����BB�Zޤ}��nI��J�
�h�d:d�G�XM:,O@��ވ��g����&g8�[U4�b�G914r�*U�(�5+Uؖ��看׼�F�;s�p�����^<�{?���K�@�&!S�L"	 :!Y�F�����PN
5P��
�~�>���+�Ǻ�:�*���ާIS�����@�m��{�)�$�9v�l�KTPڑs�E8�$84���    IDAT	Y'�V����3���5ʤ�:�����\
�_w�
�h���z%Ұ�%�a�4�#`L�: }�=�FX�<�w��Z�%$�S��.�����q�0����+��F��c���
��W��a|b2��T�����GF�שm�"���5aC_m��� b��T�"�P��;!'����Yyf�HD����Oa��~H��D$�R��P��%Z��0BQj�~�;S�B	Q&F��Dt����نjv)��뮽�}�k�}9�<�c�&��8"_*B��8K�_�}?����.�m�=(�J��,X�2RD3�-�����Bͷm��h3>��o#�݇l��@�)[���mԊ%�����H����*�J�%�!(����3��c�/OO�����}�_`�*l�D�.�Z`���$���2���2I�c�X��v
���"��E�#a.j%���|l8����q��N�_�~f��x*�	Qx�PΗP�T!�r*�k�������q&��^58՛�a�®G�������h�cól�I��!؞���C�<�������(�u��8�%k�m�+nz=�g���/�����Gss��'�7o�a�8-���q,^�}�������f�ص;�����n|���*�$�Z9$5 H� ��RT��s�hPv�����Q�nqGT�ښ�;�q��F�.Z6P�`��!��|��7��sNjl����N���j�� ��,z�aN�oooŢ�n�{�9��K<�������I��t�6����w��k�*Dׄ�yЫD�1$����U�&�D�}J�615=�X*�S��|���mX|�Z�;|���Y77�,�����w��4�E��BG z��^r���̧?���{?���顇�	D����G��Ť�� �9����I�q.M}�а����L��� �k0f?qI�A��l��+Ғ�����>W8�w��>�u�H���%HO��ϭ����IY$��s>��yb�T��s�W���ijE`#  D�<	@����7:^�����.�Ij@��r����kљ�:e���w��������������\���z����qdt�,AP5TL�ylzr/e�{a8�.Z"��KR8�/�6aba!�X(��X[ο�-/8 �9�k���la׶'p���$���@��!T*:wK�h�B�W������7�ģ{FP�#��0D
���1��Ts'fF�����Q�:��~�	+�T��T��m�i'j�e涏+�{L7�x�B�Ne�lmE�4�1�x�DS;}a3v����᜿��IxpǤ���W��\8x��t��t8���qMA��E8G��C�8��٫Z��[B��ق�ל���]�?���!k80]?���|\
+��y��*&SH���6��}9|aU��S #u�I�!�d�*.>o5>��;p��ݳ������dg/QU�k����*�H���L�����.�����Oy�d
�*#;3�+��V0&�����&��mrB;M�B'���d�$�03â�x�ҾspD�u5�K���_�|��X&��-�ɠ�8�iX��L���|�ߺu+w���k5��x)�[%DbQ����Ǐ7���0 ��.C��|�ċc�%��!w\0rҠIP�Q�7i�ȅʤ�x7���MI(�(@��D{�����/G�wqֲn|�o9�;l��}>������\;w>�h$���f�v�r�v�r����}6==�Y ��Y�ن�$��_�"*�Iڰ�\"MD�h4H�7m�&��h	��23�&2o~ǝh_��8ē;�.Z[�g���_��S��q�p?%���5W_����F~�'��O�Ģ�k�l�ÿ��<�u*� �r8���y�A�J& 4����h������Y�A�Y������"'P ����@H ��e A�`p�:��� �q��OY/#f�޹��YG��}�$� ����?? i�����\;_6D`G�����X��G��+�JX�ہ7��z�E}hn�g㢍���P/����#|������"=1����۞yƧSK�c߉i<��N���M�i	�ĥk���/��=g�Z5��ɽ�6��]_{����ѽ�����JZ.�c��S3P,��D:
�|���s.El�*|�k?����+B�L��>"�L�A(L�g�X�]�T+`�c?D�&G�3>�G�v���y��{ԅ�(Xw�u��+R�a�O,�d�!��{��T��矅ǿ�)��t�_�vO��kn}ƦsA��$M�$$�*�����]�
[�B� �̷Af�aQG����؎N�emI�O�����p�$��"�iϔ�f���b$(���8P��-��zj�"���*� ��2S(�[Sy�A�'>�.��S����f���&S�=��9��-��i�����6��K/FO��O��|LL� #�����KV�-������da���J<��s8qX�lې\��bZY�bpb���p��A�qqdhr(� �B�h�q�����x����yjF��5�W#�ˠ���C�d5�CǏ����{�g�Db�0,��sP%��q�W���4��A��Vp}H�%.ϗ�qכ���D�T�b��Rr9�U�/ŧ�85��ȑ#>�w����&Y��>�R1� �l��^��C	�i��v?#�Roo/�Tu�c��m�ѿݍdT�D�?Ӏ*�,�gG/I�I�w���=D?��p�%��ͷ�9���(�i��Z��P)���օB���RH�����	�e�-�����,_�'lپ�?�r�Z�������DY���5`Q( Q��Ѧ���,�Q�Q^{�OHh�AӀ �uMbl�C�Hs�)�sn�DC�9�"��Ȋ�S/�.�4��������I+�6����Ї�G��X�]��juW�>6���1K��������v\Ȓ��T˖,E)�Ǒ�J~ @n~94�H*��K����_���/�����'�[�~ڧL��E|��L����78T� p�%���5��~Q-�(��hWLx��I�"m��_�����߷�\�ٱ���!YaAy��C�F14��T��d�����K,�G���pl�AKA7����;���&(��*��z��xVu�
���m�F�����?}���(�@�h�:%{PU	Vn�\��}�s�ϱ/��׾ 1@ο�u� u4�:�tš���+
ؠ�sA�O!�'T8��X/f�ו��-w��5ߔCx��>����Q�UX�ʅaA�d�t^F8��swG'���$��Y�-M���a�SDt��x����k��?��D8�iC"�axx
吨
�G�q�Yg��eKR5�h�qH��h,�X<���Xq�z�o��Oh�U�:kI(w���2L��"]�y�J�"Ä������v;OA
��㣓�����>�D"�ήn<�g?۲�����ВN!��FKK��f��)<�gr��{�	��"�R�.��*���V��n�ZJԑo ��A�����OJ$8R��@!EBLn��b|�/^s�Z?�k��L��r��w>����Q�\%b16-X�n#��<����^���Q��wA'���O��>�a	*�X�t�ls�&��bt*|�z�U�i��E�Ia�Z;��7܊�^C�X@�(_j���>��F*��O�&c��F�k��(����V������܉�%�P���#��@"�H��T$��?w�=��������y`��Qb�rE�o�E��v��
��D��.,q���&4o��7αe��I�(�^���Y���ˁ��$�?�]2@�G���l� l�:�m�� �H��/Ӵ��]��i�X��\G�&{��n�;n��i����x��y �8��w�_��]��8�_���c[�-;v��(@w\l���}#�qp5!�0�.~B�q΢f�tm'����gѩِm�#@J���n{ĦU/�uV��� �-Akx��ObjtM�t��K*r�
<I���Q�H`"��F�?c�懸���ԁ*A�-�8�ŭ�@uE�[�+��/}W�ֿ{_�f�o���t��l�愹ܤO�i�`�s�����[��}�ͻ�W�x�h�u_��c��"䠫���t:�Td�\���:
	�KY�w�jl��?	&f�H,����]�{ͣhH���"�]�S�Y"K|z�v���>D5¡tJ(�x"
Y *���[u�*�U��d�|���ֆ�Op������Y�b	
9�2S��Q-h�t\u�X{湼۞x���M5���hMc��N�ç>�8M|g�3�L7����$(v�SG��)�(�~~�{��Gy��E��d�e�׾G�{�>�{gWL�
]�9�$���t>��j&6��7�e�EҰ�G ���F��%v�s�}47�M���@��"�x*�i�H�0
�MM=f%�[^u5���E�n'����㓼�l�Li������,�	OOO/V,?�'^�R�*#��qҔ��[��.l�����C�D*q���%��!�l�LLSGU/s��&Q�]�;�B\p��8<0�,��rN��B4��t߿��T	RH������k��"��U��YkW	;wm�����lzh{jJ������C�i��
\_���<Š5' ����yx@�'m��މ�r�8��϶e1��[#��)~����F<m	�DݤIMoh��ΰ[S��f�JA�:=�tk�$64&s]����YǭƋ4�`B�<Og@E �& M�$����R�`���Ȃ�$�s��ЙT`䆐
K� ���}�x_T+��F/�w90�+�{��S;w��e�%�rg��l?0K�Õ(-�@�ѱ�=���/B��;�m����mx�$��{!��}��{�xי�]~H!mD	�_��^T(�9�^5
'�)�Q0=�;>���	%ك��`<��A��0�1)�X�$��k��e�iR�D�IE��^��曰��dz�܃|�G�����G!�)df�\�����xB�m��%\�җ���}B8���}MQ��{G��n}O&t�	��e� ��v U%�<q�	(	��o�[�)���X��G�]�ّ)?�H�橸�o���� ͋(Õ}����r��$1p<r	��&H&���pDA�R�����s�C2�@S4�E���}��?}��O ��*�E@ڎBv���x�:Ԧe��+_�3V�-=��?z�8��a��W���jo�����?Tˈ)
kV8�<�:�"u�}ԥ���9v�"�ʵy���
����\(k�O8�hF6O������Ϣ\!��~>�77q�H�T�D6�'w�D��0�����$J�@,��4
��	H�+���\6�u� �0��@h�ޏ$ �zq�]���\�a�08p�/r�Uu�^�LLbz&�kC�m��r�<ѯ���p��3YP=4؏P4����E8K{�ч~��۶ ����S�e70�4�i��m0 ��E8�D�b��+�¹]�g�Mt�p�hF{8�nF6S�ￏ�G4��$)H����a�c	,���~���y����n��DV�a�a�r������P$>N�Fȶ�]�$ڻP!�MnhzA����)H*�ց�Ki�2K�"@ɶ���0��ҍ�+�B�𴳙�$�y�ـ�� �8Q�T�qy�%��IW���/4����ة�~,�G�j����̙�����0ɒ(�(�`%�1,��A)_b�*�@���[�`���p�y�>��}�y�W�O}�ȟ����
<�g�_�UQ1m���804��m9��3��t���!E��\��Kc��hkH)�	׾�v�Z�!DN����Ҡ_�L"$�����_��Ԋy$�)�t�`FQ�|�fK�?4�)]����D#�*�g
�<�J���A�K6�+˔���Ue
�/~r7.8��w���m=�_��?Gk�R�LʨPQ�kT�b�K.�j�]y>�ُ³,n�	G�-��7܎�'& 1ʁnuo9$M�p���.8�1�
��<H�(\r��mD�!��U�z�wQ,d �+�����:<�	A
��i2�j�
u�]0 !�`�|P*�$�(�,nI� �d��.�b�л��H�]��Ň�{�^y���ر�/u.�R�$&�F�m�Vha*�i����+_���fd�g@��+V�\5P�+(�hJD�z�b|�K_Dnx!IBX&`�D��σ�4�G��ʕ"J/Z���F(Մg�����::ќ�3e�0,���Mb��;Y��҄h]���ڂH4�s���a���&x�
� �H��|�p=�FPqZO����e��K��p��󧎻Pׅ-s��0ODX����X�l.Z��y�˘�O �tF����l�3ؖî`���������U�p���026����hmoAW�؎	�v8_�=�'C��]l˫҄� ��!���#��?�Q���}��cp\	gm8^q%�����ڬ�H5��&;s�9��J���C�4��#�L�����1-���6��2��o�Y�-Fplh
ٲ���	WJ8�?I�x�)ud�E��5	��uG�j|��P��E>n>(
h����X*�E�G�Ue C"�M���V�D��O5h��.hu��{D$0R�F���Q߽'5!�	$�Fx�z�ϥf��G��˓�^s�����	�!V�C�ȈBD"EOWS�Ɔ���t���7����� ��.X�����W�q�ϯ��
̯��+�{�~���Mg���-Xx�=�;�Aޔa��!Fqq��k7.��ՁX����&w扻��ڗcњ����4,�2�W�Dr���H[��Gw}�( ��X��!d+N�Č$���Pv��V1�-2��j64�@�Ѝbq�FJ4�4��(�24��̡���`�}�K�B��<]�-5�Lp3�z��
^u��������cqk���W��z�qJ
��B&хG ��j	�D��6e�K1tcI�J��%��f���'��5���l��[���	3eP)�D�tu*��IO����ap<i�"��w��v���$��k[�$FYGKST�Aw*����f���+ZON��|�I�:�F{{;jz	�6m�)����*���ZlXw�p|���1��u�R�9\�\.qEoG;���"34 U�QB�]�D��D�-  I4"��+E�x%]��j�"1���>�ڍ_=��3y�~�X�d1f�'199�Ӕ��`���~�`A��"O��>g=w�[:;��{~�_=�8���0jdg�B՚�X��Ә� �O�q !�2����x���	�8 �/Qi2壷�	��t�9���n��Vf�}�ZE�p08:�]x*2����l,Z؃��̵gctlz5���V���;Z�Qly�!< �u"j���ǣ�����Xl-M �&��A�%�DkW�x�u(�
z��b��嘘�D&�Gss+L��W��U���.Y�S�d��L��t�,Z�־7��&D�i�V��D'j	�#�O�� iGd-��U,�XgM�a�5H����VT�x
EH�v��Y� �n�@ ��i�X�5�h"��%�xЄ4<	 4-����,��Ǹ�1�Q�����P��D�u� ���y���(X��Dx�F�8ؙ,���>�cʈ�CX���4���a(��m)��nBgR�X� ��{����p��u~�W��W`����+����.r��T�W�b��3 94V�dE�-*�d�
����V/�E+�p�����!%�*`�9�j�F��v�njl���5W��u�!�a	��ñ�����f�Q��@�*�Ӱ��0��呵(�>T�4��&�5��'���g;\H�3��9hmo���	o��,ZB����Y깷����X��M���On߃D�B�O���M@��
6B���^�2|���:�.��}����5	�l𤁵����y t�=�g3�DT�p9Y[ "qt�t��9���$���{���b��L���C(ya�tz>>�s
2��N-����e]9��˪�nDt-v́Ov�>�+�F�p�M/�矉�d�C���    IDATuk��m߾�X�U��b�������Y���_��/�06>��߻�"z}��%t�4G�����ˈ��B�~ @Xe\?^��0�E�2Q&��P��V��=�c��_=��'Fx"��wF�155��E}8�?���x��:;;131��}^|;c�]�w~��8p��MͨU=H
��&x�A �>�aaOn4���� 8�N�w6O l�*���N�&�PYz�I���.O��7���L����&ff0:2�t>;�y*�,D���W3h<)r�D�������ґ~��b��Q����S�$#����2�/�*;  �u�}J��Ś�J�{���CS<\��L���r�i=�ju�=���e}X�|9��i�����Ԅ���02:�7�~;��yR��"o���h=���i��w��ę��#������'��ȩM��J�ٞ�X�.d���o�OA)\��3րQPg�L
��U*(\��Ac�b� M&��(�7�3<����t5Z�s�_���?�#���f�Qz:���� i��IMI�~��NS�&xB�ՉH;��W�@���=�{�x=6kp��<�`ü�|1����)���/>���x1��Om�mׂ�i;G'�x��=��� UӃ��ݽô����Ugvᴔi�}iaɆ�0e�}��j�h�[A��o]s�l��:5x�	�2��@�\�
�x��G`V
�M̓�˨�
~���0t1����!�08Q��L ��
lK	�4�@4+��iO~b�������^��7.�����X�_��"<ux����G��o���i� 0��p"T
x�W㛟y�pll�_��&�=6����D�
a�� ��'D�
���naA�K<F��yB)��p��\xs�X��_���012���.�п�ßžcS�[
9�nf�A%��@�^6��<u���"X���!n�sad�U����^�*$�CsD�?���p��/�u�'���p'��7Ń'N���(K�_�,^��������h����3	T�CW*��}�����0����T��Mnh�@ֶ���� �j�0���K����"�N�/U��_�eY���3IA�j�'�D�P@4aJ��e��׻�J	W^}n��&d��Z�G8����G����!�Ʒ��*�� $0br9h��2O ���Ё�'�A��ZH�����jcp��S�㖧��Ŋ�:���0<<�"���/��i+Vbbr=P6�0�.��Gaf?��>ȶ���!ED�c�d*�i�aԘ�E�f݆I�Tsp��Ţ+0��9�)�c����.9V��Ol�¾�hio�)G��V{K;��:���?��k6�p�x+�e��Mi�"�@�����0:9��cG!(4m��eIc�
�U
�d�\�d�ޠH5hYt�fACC�CZ���t�o�	9)ToL"fKT,*��4� (/؍[�Xc������u��Ӧf�䞜ϡxq��d#a��꾼<�W�i@�$��tv#�ɲC\D��W�W��;b�N�@s\�y�7��>�_����4����x�P+=�:4+���-�'	(6-��cy���]� KC�� �r ��~��:n8�4���bIZBJu`�r�]��&�-Z�u�_-A���dF��F��ϵ�e�!x�<ڋ�#��/���-�T�£O�Cُ�y�Qq#828�2�\H�P	�Ph����H06�l��dH�׿�y\w~0�922�X�@�,�?��&����p��S>OM�o{/��؏Hs�ܑd����ùk����p�cn�����?��Xj%�F�!�p�@�JE��� �ڰ�p�E��Q������^v�:|�#�a��at��㬅M�͟�W�7��hG�
�pm�]��;�(�V�D�-�p�4SǏ�R tw<�j���V�BU=DU@�u|��?�׽ꥳ���=~�X@E���L.V�`�[%S������q��;���=5ӄO�E@g[a�����o� � �0�i\�tkݕ)�PO�]�,�m�rmHRq<�s�Ÿ�+Q�=�L�[�pitzQ(W01���C������]ҷmm-hiiC�\�%W\�[�x3�=1�i �fоQ��B�4L�:�vX�0B��֑�n��(>�,@���kN�CX���&D������]�>�<�W��3A?J�,���@Z�ZY�N.M]�<�(WK�~���ʮh����?�	Қ�w!�.�)��!��,��˷]��v,�AeM�A@41\���t/Y��^A�61��A&��H�+����MNCO6őHř�G���֕H$�q��?�������0�H3��Nd
l��"%�ph]�0R�� �,
�,�j� ��Ҳ���p�%�K�\�d���pP{^j�X�6�טt8��,�����lB�������\����I*�s��������j���uk����'O��^O�����?"i@�XԵ�C,'�Ǡ�>�b2��/ބ%�q��$��?����}�@_l+0����������S;�����-����=�,�O��*2�ᱽ��oͯ \����9��q��%�U�WF<"!WȣuA/V�Y�ޕ� BBt��u�Uf���^|�]�D"���L�ؑ�`�;ub=A�Iŉ�������(�b�ֆ�!���aXn��W���O�%��X���T`�Jp�n�����+s�1͔���} ����q�o�_�����#"4B��D��Ǿ����A��5���Y�+Z&��*�����spz��mkzvؿ���\������$�<[D˪��o�ox�+qN_X8����5��/>�1uBQ�"��t>��7�<3�b���i�ֿ�����=�CI7��U��s1FnvآB����� y
����Wa��~L��BY��rQ�@��!	��ɫN���{��7�8�^�\>�M�|���#G�Bt�z�!D�jok����Gǰj�i�m/r<�Y�|)�Sc����(�r{6\��=�H3��
,�`Ѥ@U$�ӕ�e���d���u�q����
���n��p�I4���V`*����$��?ӱ��ji�"��6s�LʹqٕW�]�� ����F�	�u�bz�ߕن7�nP?�t3�A@��L�X��'H�&w&���4�R(�4.��ס�@[B��M҉�A߬���E>΁�8t����-����h���I>l�YC"���E(���/~��#�|������h�x�$�&�9M?ꀝ,���Do���)�+^�:�/����|EB�R��v!z�X�u��b�(���tut�{���%��'?����G�P�iBw�
�La�./'ِD#��� S�Tx�K��u<� ���0�do��MnNf�\-E@�#��I �v���瀃�ֹ�F�v�TXBt�ƔeVD�\�<��Jz�F� �����$�W���|���}'�%�Jt.I���̥�G�X�p���0T�;eB $U�)X������Ǽ�W���F�}~��+�$��E�s@�P
�:~��m80\@E����HT�kB�u��^{�z,R+�ƐV�)͆c��%5�.�J�"�A�.���{�uX��Z�G�*|�I�nlJX���`��a殓M,	�!�`�1���1�1�v�Hi�R��"C��c��P��S�$J��^�s�ͫ��.ڀw���x��˄݃�~"�Ē�&|�Ǐ����P�-D5���j|��w�{���a��cS�g��U���p�0Uꔂ�Nk�K�r�p<����>{�~l�K|W�����C����Uƣ����h�]����_���#kJ���¨᪋���?p+¾״�	>��_��=��h�<��:S��O����7 1z=!���-�W���}�0=<��&ɨ�<�a{&��f��[�;ߎ3�.@D��Ҝ@�Z���ӆ^3���.ek��,R�=#R�������*�H���L�)��iK{qd�x����Bpmؖ�h4�H$��)J�'�Ft���NX�v�*.[�?���������݈,G�,�0��::�C��Q5L���`��eL�"Z�rp��[nžバ�0j��֎E/0���p`0�N�A� �pS^	I�ْ�I B�`ʕ`
H(߄r2T��<�������B/d�W�D��0m�G�d�����3;v�\*0�J�<a8�%���!�|4��8���@�D� {^ �B�@R׳؞ͩ�$ɮ�~�JE�a�kZɖ\��W�u�L
H�4�4J7�ry�ed's,6�'chik�Vй��i�T������Ï<�����f�8}frULM��2LP4�j��X��BSL-I��|U�E�M����'�%�57P�\-HxD޳��u 2�35�P5��K_��$�n�R	.M���-g)X<	���: �=� $�,�<�9��9/>���k���M�k��@&Д�M �0��$�����|�M@Z����۰�%�jf鰌K/�����~���o~��� d~O̯��812���q*�N�Pj��]��`�@���'i��p%����EJ�pβN�Ѯ@3'�D]qa+����h�-��\�E�VR�_̕j��YߺDi � ���ˤ.�Yr	+@4�9��4~��=�;�Ū�C	̔=�92�]D�&C�t���>���X�I	�W��lJ'kQ�5PУdg�^����qú�Y��D�o�hƓ;�w݃�;�㴕�1>tɘ����x�k.G1S�Y�i~�ֱ��ƿ� ��bM0M�c����_��/T|J�^��]�����S�^��f"�����
��q|���UrP%�ښ���.l��v�J���1\�a-��;P�.`M{Z�?]����ă?/ԂP"M��p(خFT'�Awg�/� @�A,�Y��`�ow�4:��^$*dGXǭ��*��!kX�l(��T� ���h�vaXf�I |�J	U��D"��.���O�6:4���z-d ��َ��l�qٳaQ�S�@�N�& E:r�"Q1�\�B�$�*E)�����t{'n{�;x�?:�p4��Tz�����}��qbd��/�N��G"��j�^�ӗ,.��:���0j�����#C3��h[���W�]=���T�d�N�R�I�^���S'Aǝ��lRiBb@M�����êVɒ�a�����=�KU�?��NL��p��R��q�F$�Qx�$@�T��f2x䗛�
l�K`SA�OB���橨�����b�׆��ga��<�_��5k��ىP,���C����L��1��X��hQ�dCC'x� �뮻��c�01�Ek��v���?>��0M�jDOTT@V��CױiA�F �[H�/�`"� ��� ���` P/��$��%�3��O怂��# MF=��B�w�X���Ö7����N <��� ��	�I 2��s����� 8�V�	�q;��Ԉ��>��q����V�`bl�' Mqx��X���FRq���6����
�WW`��WWn�q�+00<�OP~��"S��T��~��]Le�P���㑨��i�D|�Q���$��5#)���X���W����Ԕ���%�M�����zг����ZM�����j\Ÿ�MA|�3'p���� ��bll��)�$�9,�2�-_D�02U�d�A���Ơ{Q�RŪ��"JU��#(a����	�n9��>$��\�K.<w��(g]�t�x�00^�Nu9U�!��0*Y(^��'<�)2�#�J�7;��O~5W�d��j�8cA��mH'#�G�N���x��F�2�*�i�_��YE��S䑥�#�����C��$:�x���lt�C���?3_��ք�o��ǚ�x��=(>TJ�7�ܡ�a�*��� (*��L���#�bh`��l�;UѸ	f�)B�y+/�%眉���jI �#V�-dQ*W�CN:����cht�O�N���_�Ӗ-�m��K�D�r�Xws��~�t8���U(峐KQȎ��l#�� 9<��a[�PN��@TC���7�v#�ځəi��6�@�>z�����Qd39��I�z�-�B�]s�e����6N�O`|*I�bQ�i�?<Q�B� B���ȳ"a�D���A�\$�]�c�vPi�LRJSq��8*HI�N� ��Na�GX��޿���"Q9��qlؾ�l��A�B����;�6�r�OM@Q%�LN �N�`��8w�X5����m(�KLc#q>��\���>%BY��'��t���+W�djib>��F�����B�v:W��Hh.�E1\\}�UH&�X�����@�m���������gQ.����5g��u.����fAU"0]6�:YArA/L��?B�A5]��vE�ct}�' l�5��X4��g�25D]�O II��-��͡�&^��렲�U�l ���?<�н���R!�&�A����LD��E�z6���ÃO�&2�`��fs2���f�*�&�!�E2��o����⚀�7�k@�$��7�Y�y �Y���cY��'��L��u0S��d�pCMx�7{���a=��Ω�T�S�T&.�SEL�a��4V�4�'��ގ����d$�^P���p)�s��MM�"a������
BT Xz���J���e�6��N!q�� *a�Z��Ǳ�i���L~�5/S�#[p1:�G�R���`Bt��� U k4E���ӆ��X�Bi����8l����c�b���(Atl�À�g�}�����������׿���VD���^�☐ky�?c	>���%C��銿�-&ϛ>ѼN�=�/-
'J>�ͲX��L�<�������~�	߾���b�0|�vMa|��H��g�[��J�!��
P��ear�u�����$&��G��c����܌ǆ0�����FY�M��$E��R�����6���W�9���3�R)ϖ�OMT(J=�0���PQ��ݍ����ŋzA�cD�!PD�T*�az�ǏíUWT�wԁ'�D{�����X�O��:�����t�R���v�eWbɊ��x�$�$�4,<��gH�Z�h�RNn'k��O[�2o��ݏə,��я0�/�j��m	��bjh
P"�CI8�����bS��BQ"� ���& ,<�'k��l @
����dK�]�k��hkmb��Ζ8*�O"�:�05�a�B7���2�4 �����!<�m"�B/
�BO�mX1� ���ٶݰ`9N�0V¤���#�Ɣ0ϩ��=��>$Q������#��?�V��E �r-~�$��B�Z(@���&�q�S�8���|��\��V�����16>�vä�`d�jH�,�'KpD�����tR�M�� /�ӿi����<5����$"�4#4���E<?ƍ���B�S� 룮�ӷ�&���	.U�o�`"6���ꔱ��� dvj�v��q�9�F�?����{e����9�OD{s��ML���L�3Z\�|ǭX� 	#;����.����X����E��ϋ�����
�9����]�L�EM����[���!��N��L��2ǪRHN[�8���I����d�DD����E��P$R݋_��,�3>��n!�HxK|y�D%*�T�д����+�8:�E�Q�<���D��2�*<��Pז9�.��A�B�IA�(��̢X��Ã�~�M@f�t,a<�����O�P�a	
$M�˚��C�j��,���a�����p�U��Vb�0��e�A�s!�5�d�Z���+�ne/lJ&�,�l��|����$�O��@)��ɰ��h�?�����a&_fmN�&�� M�`�&�}V-���#J
5H6���X�Q�Ը��(i�-�]�"aD��HDz�tc|��ŖǶ!�)"I���B�F .,Su�e���5�p�X�ь���3��G��E�|��U��ƙ�E�崷w���	-������`���4��,T�UI�k�� ǲ� �h7�"1B��)�    IDAT�ܐl��E�-m������K��43����	ȡ(Z;���g���Z�x mmm|i��8�r���Q��B1n��.d2DMC"��aB"jМ�k��P�   �C ~}���9r���{>$Y�L:%ˀ$԰ti/��x6oބ��c��#!���Ҵ=v�d��U��X�믿G��t?�Z�mm��@u�c�{� � �	�[���@CA�q�����!P&P8��,Q�9���M�ri�8�� �� �L�r �:�v:��ή<-�)�*S�BC�R����fq{{�t/���}�`X6OS�Y���H-�C(g�Q�c�A�/��y`-ȩ��d��U]�A���ѯk3(��<����������ȶ��)`s��:��$ w������,�1ڨ�� ���&ެX����S�h~J�4��6B	� ���	M�4J�"��v^�	�%�1�3C@^za`�=�_����W`�����l��+�s��P�2�Aw=��dL��|����t�h6$j-��O�K��L���z�SX�"bu��:�V��_Ê��$�Yb��0���>JצoL���=��{��L� s�55�_��p����c�TC�bat���)����$J�
�	��P5�^��gDPAAJT�=���Y�C�9���6���o��~�Zlڎ��/�?�EQ@�p���PG�+Y�E�"x����W�E$/�����`��4j%�X��u	��%�[�����p�ek�y��K�����[�I���p�������߄��i$�ZQ�-��VU������Q|�}o�+�9!��S�x�u�]Gb.>�\S�ar����M\�`R�Զgq`�<��c;1
Y	�e1�Iv�q��T��,���(LO0v��P�rև(+0,��a���Q�B<#�[�֑΃@���gvXr,N��"G&�J����	8QB8�<�r|�ms-[g[e*
IcA"x��$Ҧ�PGk;�,��A�S
z�VÉ�QN�^�z5�߻�;�*�s�"��E�(�6�P��0>�������"6[r���a @HӞ���#~@��H��;��I�3��y,,a����Y�?��}ЋӐ$2Q�W�f��*��j��6���126�gwl���s�D���d�� ���d5�Z�A�M-d6L"�����gS@�]��>*�x�+�9'�s@�"m�z��w}r��h��"K��:+�� �6�Z5Q����ځ�'9ٜ(E&k; ��A����K5Jh�h�I��3@p���t4�A�`�~4٫�'8���gd�]�p�^��E �D�R35�N۪��_��[]KB ��'���!�j5���1'5 ��,��M��q���A ��|:r Py��F_b �H0��N�$O�CYnz
!EB:"�}�|#�u�n�{����O��k/�
�_</���?��
�ؽ����T��B�%���'px� WN0��7,�"y�ȁk+��pI0�XH�U�'%\�nR��:�0�ֈ���ɭB�MD�P�_�E�<�&�Od�-}aҗ29�P��:�-q�E�ja2_E�j�P�~B�	�E�P��860��QE�V�C2"���x<u��F4���}�4�I&O|��˷���7��M޵�������TOG�"���D�I��z�g�_����]hkSq��[�~����&P��e����{�sdDF�sVf�EM"C��P[@P�Bm�ѷ�[o���j��n]ح���-�,�"
XT�LMԐ��<gF�|�����7nf�"U�padEܸ���L���= 3HGP].#�N!Ě�TV������ލ���wC�Fʿ��R�u��60?���=�'/�8>�N7�f��t�����Q(��=���-oz=nڻ�:m����ܰ�#����V��z�iC���>v���A���>�5kq��1����y��W*�@�h$H���;7cӆi�?}�~��lHuʣYo���dr�b�e�ڤh�J�ga���{l�pb�E]�QaXĵc��[�I�n`jjR��u.�ϡv� ���Q"�w���
9�:w�k�q���ٟ�N������1�U`����
+��(�^��D����r�,Y���m��;ئ���5��$�U{W˚3�,N�<07�HR�y�Y:axd�b^�\�T9�+e�=)��3���@�'O��J�����%�C�iS�����ӎ�_��޳���_��yP�f@���	�'g@�+�����?� 0m׏ke��笊z�����+r9��TA�"��f�`Q�&�&=�	L�;�B��O n��//
�	�M��ݣ�gy!��TEJ"�O�~�<�7��8jW�N�a������r��9N2NY�M�K�m��u��}Nk�Wr��<� �T� � D"xyXZ;���	5{�SA>�-5 �`UVL�K/������7�#�-��u�-�j���3~���9+0�x�s��`K�V��g�s��H�2h$��!���>��#x��94�C��@�$�,���[�e]Y��Z���͓y�1TP�H��l�`8J`$�09�G����N��
��T���g� ��]C��j������*�$*]
�I�ʢԊP�1_jb~��J�.-YS��$I�a�jX|W4�A���M[�\k��l!��o(����D�(�U�������Iٸ���Ni�ј����(//�U���O�.��$����?���#���l:)-���ȧٱ%�,)�RvnY����)fQ E���#���`#��*���,DI,/."nV��������D�SL�m>&x�<��p#]+���2�t���
���2Ry:*���8��;r�*d��h6H{kh-9Uaa�IA��{�h�mM9��Z�@49YLXOe2V@�TqnS�*��� ��ާ�c���~C݅�/$�u ����:�d�`�p�E*Q��!Ki��^7�0� �8�4Ҵ����RRQ�#�#v�	H��w����Og@�F7,��|���V|���!�)��n:8%2L��xv�����Hf(g)�H�j���@�����Μr�L��:�>��@Er@�P���#I(�dq�Kt��&ڶ�����pB��¹<itI�����M�bW�k=�� X`"r:v�RPA:�kAX��y6��捨��c�}�l
b���*7R�D�} �OD���ŝV�qۉ����$�&5�'��x�ܑ�[�M!��H9>�z���w��q4�#����&F'��aב� V@��r������ ���\�b�]��Ţ����9.�(�0�X?Y�Ͻ��6SDwyVlw�z렆�xn6�������y�[�O����/�/"��LX�7q���'��$���	�b
���k<��w�X�7[�&���F�j�7\���*�X7�ƺ��q��Y��:2q�C)���$�5MRh�+�&w���ڨ6�Yf�B��6ʍ�0��@��r3���u,�c����6�9���T`�If���	�����X��0�B^�Vicԭ��ʮ���
���.KRrDHbױ^E&�E�N��ܻX��HR �E'��e(y�)�\�j	A6k�zeYE|����;Uǒ� �p�0�4��Y�TA2�����N�AjdLE�N�T� <`�W�T��Dً�%*�
���|��<y���������9k�K�<�Nő���z��t��W�ZU�eL/��
����/�lBa]u�G����
�ީN��(�I�����$fv]\�W����tLk�TP��	Z�T"$F�[`����!f':�AF����V��V���tG>/%H!��Ȭ�8Y��$�ғs�r�p{�-����l���ΞUs'r�N�OD�r�,�2�H�j��Y����X%e���	��n-�ad�C��c@�Y<�X4�6uid9�TL6w7��l�d��#uu��nVڏ�o\-Ԃq�G�]̉*�A{����y��Ϡ&���s����F~�fTh��I�������ߒW(K(7e���m���+�D�lǇ M*;nL���FU��i����)���TS7�"�=�I������%(U"`O�sO���zᤋ:541�fh�w,�HĻt阈>��犻�x �sgrl�ffP^,�̩��`�����ֵtKW�\�릛5�?ѳx�/�\</�c<�ÿ�
>q&�0{�Āb�z�������ы��mԻH���2i���%Y4��Nq�t*�Vua��b����[׎ar8BЩ#��#�)#Ѧ�j�$�*�����z�Xvb��k-ĩ,��"I1wT�R��6҈�KM\�RRbr��"��u�:��J0&\jP���=���LL�å�y2,()��٨��Ҩ�����0n9k�~ 犥z�5(/."��,!�:)��h5!!4�à@Yq�]�ѷ�@���H��
RiZ��[cG�"�����H�ZYYA�8"�<?������G�V݈��l�T�_Օ�p�p��椁�X�KX.'�-��`�[*�ҹ��ͶhS�\Z���r
ETke��w�q���z��fg<�}K)-�(S�?������"�z�'pbE%ZE�I�Ľ܏���/,5=`q�w)�:	Hɡ���t1� ����.QYZAyyEq�#?<~�4�q��,�5����
K�K�N�5p! ҟ��>|�^ Ĺ-�@(]�4�s�s�I�� R�G�ᱦp�|S�X��E��\`�>MY�$��d�55}bC��C^ל*q�d-K�:��T��$h3k�w���j,���������4�9�z�(w�<����|p��ׄ�k�z1�bٹe6m@��FH�c�	�x�px_��M��c�1�o`49s�r^�l"(?Dѐ��y��\�k�D��1���k2�th|��U1�ޮ���6��e2�t3A��<��ŵ7 �]�cjܥ�:w|u8��L������9���c�Ҫ�8vT.X3�y��^��$��%q��
����:x�`�Z� ���[�g/�g/΢ՎQ��v�/-�����shE4j�-$�dB)�MO���y���ޤCTf���x>�5�y��0:�B&dxݒ���(ZF����MX�&�F�f��"j�$��.mR�F�Ri�Tibn����
ZTO#T���j�e�Ү�D̒h5�v�N���D���y+ZX`�`"����ui��@g��Ĝ�¡s�L.�O.6�"N��'9��ј��;�윪@$-�p��N�M������|Q\xN=�W"�x� G����(��E[��ͪX�N�\��s�	��I9��?qAhb��6�u�z�9r��9�Ǩ��6�)�4e�ڲe��f��0��E-�ν�{F���|X�d�o��x:�h��&�N���V���!����`7��:f��X�W6��VpH18�FT(H+B�0:4�n���+�H%���H�Rp��U8� ���۵.���=YV����$���q�P�<�l�:�S�\�s
����4L��hm���3X%��i��+��IV�m���L�ς�t'(��<_=��_8�4�M4q�,|�d��q�ݓ��n�H��qt���P����,��Z��� �� ץ�@&�����8{�Z�:���߂�Ĺ�Z}�;L� �.k�3TP��tH��t��H	��Q�z4:.�]K$P��^�M:����
���:n�B9L	(�39�V0::��
]׌�) ��̷�s���������#�n�P�G����;ϛ�B[6o�ԉ�(d#LE�ş}�&  4y�wj�A1X���
.�����셹��_�/^YP�W���I���%|����w�lm;�Z����;��p5C�p��$�o�!$0�Ka���h�)�5�3��(�T����b9��[���Fk�&���hw	F���B�j�Z�jC A�Ŕ�F���=�na�EzC��]��]$5���42n4'�]�-�]`Oh %�RMX����x_�9�γ4�����O�L
�F�:���\{T,��$7��7�E�A&�b�4/��Ş�cE�/Y��O��-�"���Wb����Z];���N[ԓ�6�ԁ�h�J��x,4:%b������4VVV�>��S��i�֥��A��i�zB�.;ɚ���D��4*���ERS�n�ʐ2�S�4y��{-��-i���p�� ���X�N��ф����0dR��SG�ͪ��	���,�X��xu�}�\�?fV�~��z�<\Qj�w-ɔ�^�s�V�̓(א.��#'���g�ٹ�.7�G�S���T�E��-��4)f�c��`���5VxKS��8���߽����51�8���SW�� ��i��&5�b��N@�8>�xtm�W	�3Qg箠C718=5a^�毗~ bֽԈtDٓ0����5�F4�5C=ϼ �PQr�g���;F��ύ7g�$鬉�F��l5E1��)_�#ٍѬב�B�AK+e��ע���U������ ~Ŏ�ճ�u�����]$K�$P�f�m�V,�-����_S����^l��#Y[�+��A���շc �۱ʃ�xެ )X����`����g=�g�^�R���Iҏ�t"���_�x��
BN������ݐ@�EmĎ6��ҝSaW�&`gi��bK�XahZ�v�lUS& �� ��*��PvU���E�s�-lp��4R�����9�Q��C�;��=�����TdsPѕ�ܘ�ذ@	��kS�D�,V<�D��7$]��ALZLB���[�^P�.":���IaAAqv&����Q�⮾�Kn�#Ȣ[P���, �{p�sH`�*o	j/r�CML`�}�6�1v�߀cO?�V��v��`;=�NKT0�V۶3ҁ����* ��'��,}�*���4,���YJ�	q��d�`��,�R͙I_
T3{Q�5 ,�DAY͘a��4��Et�0�G��d�l�1w�"��5t�NP�o��:�Yȧl�����
pO�r�ds�k �6�M�����]��Y��٢��S�#�ˡᜫ̕��,|ٱo�@�
~����pZ "u>2M�zay�`v��D�vq���o����A}9?��`�ܜhsK{_�1��;�����Q�.ϵ�&�7|Q��h����&�\�t��I�>hQ%���tk�z]k׍��y��t�"��!S,X;sih8A R��t�fY}+ b�l ���S���u�k�07��xO�-^!36�L��x�"�D��?�uM���9��e�@h}�Ϥ�c�vM@�9�".������Il��!��:����6���|��
<�
 ����@�
<�Ծx~aA�A2�<�,�<~�}�����z�N���W�.����F*F�д
��U#FZ���fG��t�6K�9�z��02+�Y�u�`���R�r���H�Y~Q����%}��)��>��9�`��-axd�������S��c������uYC�	YqK�M����	�X��;m$i��ZA�����VWQ�%3[�b�	�	�5Q��d������	H�����	��g�d�;��)� ���N{�AJ�M X��ؔ߿
~��Y>CB��2DIZr�F��3$�����q쉧�\YF^�XM��q]�$]˜��QѴ��V�nA]^xJtf*�$<wT :1���pH�CA�M�8�`��$����j� 9��_������2' ����I��Pbu�';n��qe<�l�4�Bw���,>ۏ+����wL�,~�(�2�W'��Z�k��9�����ti���V�BL+`N�Hws�P�F��So�m�$��&8:���<O)�F�h>�ې��Ӽ��w.X&V)X��,g�]��}���Jd퀁L��h�L����c�F�I�845դ����b��R�I�4�*�＞����d��	��!R�1�$0ZB�\:z(�Z#��$�X��	�y���i���蚳/^#�q�A cS@�{��fg5���' ���5�(��	�����6��N��*���O@z�z�߸�.�UB�K��H d�Ν��>�?r�U�Mk� C�wD��a�� �������n    IDAT����_z䱸T�"��1�]w�8t~�{d?�_B��� �����Y |u��UT�8ЎB#:�q�Stni�bT6��.�4J���0}�Y�r��n;�r��n� mG0ؖ���6����k4Dnx��G��z�	֡U���N��X��+j��ֿFV�ΑG�r~ѩ��:�>��5J~v:ɹf��$i�f3�ЪԐa�D"�ҥ+���`�B�LM`��x%ē�ώ�e����8�6"����U� ;�l���uEU��3��H�J�Zض~N>�O�`�oE�M����o��@�J*��{wX:���~�w�����ɬX�w2�B`�+�\a�B��z:��ȢpT'����`@�P�(��'uez|A�+�����t	�h�+T�/��A���	�Uл鋷�u��:ώ�/p��ZM�U7�>P"a���u�B���xnי3gD�Q��Q��M�96�F��Rj��é�@���9�[���4�U�`m��4bE�(��V'+v<8��E`�����:)����/�&s<�(�=E��
m���C<<d�B�t���_}���a�M �	��!�Y��t)ЗVA}F1c�����.0�L����%1�vZ�h$u�& :ݔ�MBlķ��m&a��8D�T�z������㘞W癧���M�݋�R�D�(��m���g��,*���|������)'Hb�= �=�b&��o}�& ����� �����>}�V` @�mK=����
<��S��JE��D:��p|v_�w
�<~����N���*8�l.����U��FC�+�wȪ7f�5�XM���tڽn�� �Vl��u�UP�����*��0%'_T'���'�1:>%G���y��S�. �
,�6X�{�t�G���8���Z�hJ���\a�J{��Uѩuwٙ��R�f2�K��h���%S(��[�<k�\k7o���9�JKٰ�|D �rK�#��'�q������a�	[=@7]��a��M�kq�}@��x��, �@�l?��vN^K��k����;���� ����{w�Uq�h��a��)K�����߻Iw��K��BL��V2Ć�$Z�<tH�sE���4ҳ�����FH�m
ٹ���%`��~u����~��5G��eq���������붻[�U(�����4�,8�(���<���&JK`���IA2�(�U*���PSNƤKq.[mmN���]'m/�w\d��6P�Q}���n�Yʻ�1�����َ�"1:" �iXÃo
�ɛ�0ܞn�q=%��z"�8a9'E4Z�;'7|�p?ل�u��|�(CÈ��LM���n�S��1#<wO���`�s����rw���}�2\�(��,��~�,&�l��PQ ��'��������˘�_D6O���i�� Ϛ��^
Ҧy�����\� )-����D!��N@@��Ӹ�ƛ5����>����\<ߑ�e�Q�\+�������"�݄�Ɨj��[�W��cG�49� ���^���g�	-	:���F�K>��y5�����mw���h8*DdE����m,�@eQH�2	v������2{�_L�f���uarC��X^)�.MG�6�:B�C�����{�G�q�k�VCG-������rX�b��b�!��,�	,⨓��l)�<F�-��U���OZZ�c�u�p��qǇg���y19�n�)4�| q��W�ML�ww)�����E�l��Ʃ��]^�D��(ڼ�0e}M��ܕ�3���}7{�	휢8��K$�.߁�b^獳NUq�/w.�MBT�9���gk뀥� u�ie��*�.�k&�hmܯ��ku~�ط�M9l��%�}���M�A���MoԐ��x �>�?~�iX:��}� ��x�|��i_�N��>�Ff�V>\r��Y���Y���Q'y��偟��y`�)gv�آۘ����"�oԺ���<_$����i$V��ۃ5��z:��K4g��!E�r�s xdI��:��(��Ϲm��'m��Y��7@�d��*�9��,e.x�gj�xk���HV����dB@�����pϫ_�O��'5ya�����7��� ��A�@�ϲG�ƘY;�\:���>���(&F�QY^�����l؀�{����c8z�8R��N�%ų�cW��y�kŝz�y��:�9=���H!�=�]���%��)M@�G���H�^Y�X!ċo�mPC�s=����_����?����\�c��ŗ��3W�$�To��\�=����C��G�)Ü�x���F���XGnW���!�G�ץ��=E��5H.G�6z�oۿ>���/jY���L<�<
�UL���ԖMh��j����'?,�m����6��P��
B+��<����b�ޓ�� ��X�7>���*�{2�P.�-7af|���|�h�޺���7!3T�o���f�h7Mxjuy��L���z�*>�?���J����Q��Rl�M�p��qT/]vY
F�Q���WT`��ka�a���ӡ9��9!��M�zˣ)'iV<�w<��a<n�������$5"N{�n����t�x�l�ᝩ��I���QXC"�/���3��������.�ӔP�yC� ��|����W���L�$æN����X��]=:�iN�x�������o:�9
�U����t>s�l�-�ג#��N3�-%�6M��N)�rK��A�gI���`�޽�DtK��'���⢁kN3�9mp����ϝ���u����e����&�������t)�P�M]M����Bݡ�4 `BSI�z���^�#�t/����W���k<��wN@xo`M,f��nj3�����ɐ����y;.�^�_��Y�t��޽�t>g `�?�$��p�'�j�x�u�����064�s�O����(/.`�M7����o<�ǿ�$F�F��\ұ/��*��I��	��y��j?Md/cj��F��������8~�0Ɗy�`��-�Ǯ��JBϧ:�̇�ཾ�V` @���`�����D\���<)5�(�b\.�����PK	�H���<��V&��|��ߩ�䗳�U1+?|��ea)[W��'͢U�|�����f��H��ڍ�=W첓�a�����%�*PE�U'��.7?����|�n,��Գ]e��~�
��� ��GO$lp�-���_ Ad�U��N�s�1Ǫ���ܹ�6���Gm����cq~���W�06���ǁ#��a�(|��S[�U꒟�p�|7�O�VS����E��G��|�23�+��a�Ҭ���}v�&N��:�}�ţ���ĭka��!{)߫R�z�8Q����p�ALb|��ِ^M���G�'T�?SF׮E���*�qhfQ7��C�4[���T$���d����_���;�U<zP�0;<]Kۦ\�� �ר�G>[�Y
�@�hM;�o�rQ�s3�}�	�y*�i�P�A�8:M� �r��)���a��W�C��8q�=ݮ(<�Z]�YlW*K:w)�:�]�r�#3Ӂ�^(��0��t�2����4�H�H��"�F��E,Q��������	�?��qTHb8��]�j^���Q��Q|����׾�5���1�fR��ԙ�:��;%�_��q���_�Ȃ!R��o40��l4����s�6�,-���C���(��ĺ�����j�� ^6[�{U�!��lve��'�a���ڑ����&&ưg�n\<w'���p������l�@g� � ��J�{�� ���z^�_���9%�sh�\��b+���x��eT`9 �s��
��& n�\��t/^%/=�00�z�.7�����B�~.�u�]g':��%�|����J(% ��e-z�f�0ZD��D"��8�LJ�{��:DQ�r�e��E���D���q��N��7~����m�k��t.�F�f|tZ�&lݸ	�6l����;�ML�܅8{邶����I�S0���������a���(L"�ja$����Ԗ����%'�b�-���U���+|-�Q�: \�U�z�M4L ����5_Za�:51*�xs�~_<�7}�t�MtjF)���B������.f��j�N�ۇ\��f�f�E�v�8w(&���^�j��@��=���O�m�[��I�t^;��I=
�����XP��Mu	��:��k' ��G�����������[���+�#��Kn
��du�& R��g��P�z:�\��!��(q� ';R��RV�wL\�5*'#�~��V�i&�R������ ���θBCT�fw}�������߬j�B0�}g�y7\�\��}�ILS����h& iҟ̥��\5
�kh,���I�Z��h��3�th6��r(r���RC�TBynQ��iMK�"iͨ[a։/q������^���<gZLN�a�����9x@ ����u ��c��h@���w��
�M+0  �
~�]�O=W-4�-���4�-��?����R.���S��^|�5 n�T��I�4�ې ���)B��Վ�N��;��9J��XѣBf*q�*>��
&�3��aQĎ|��qM?8(��,9�d���'�C50���?�����5Iw	��b�5� *FU@[�����l�z�n���_�V�Y�`����zCy�Z�kP�TQ�՝u.;�.�N�ks��Bm��U���i��}����uZU4�mU ���n�a:;ŝ���T�*RxLb�)�)��L����ގ�Q@���A``҉ýG�I{c�*w3�I��j����%; f����܄\k6�G�j�D�����uҀ{�)s3����Y�&x.*h=t]{�Q(�I��z�ˏ�x2: �e�v��#������ ��W	̳k���v�J�F/FvS;�����l���ixW-�L0�*�;qڣ�6���(ޖ^��5�	LtN�>)X�ذ{oz^��LI"���nwZ�j7FX^�(v�2v��	4Y�s��a��͘��G�ђ֢�� ��@�6Ix�qTJ'�^ ��D���y
����Q���n�NZ�.�����É�P_��d*ҚR|���/Fu[�:� ��� ��2	����l���v���V�]>?�)�"un���S��:��ЦV\OHݟ�M�N��6�-��Cعm;f/�
�L�a$����ďb��Ii@�F2��5�wU�0���\<���9x���
=!�]X@��D'�d���|噓���Sh�E4�Iq��|Ňq �ٺ���Vg��Ɉ]>�z(D'h ��e@܃XTg�ɗ�SUb'B'�P��� (�U!�Nj��B�N�v��%���{�R*�M�i����/"�K��Q��V�j��B��0^5�_�D��W�l:c]OR�����"�5[P��qeA�P�T��O�L�����.VZ_��pbc��_��Q/l3�3��]Q�;{��މ.2L��м�@ci  i������P�kE��꘥(9�.K��l�����}sO�`Ւ�6���U��.�H����г�0d�����`!���c��-ht:hvڨV�ظq#�A���G�F���պ�<�5	ӹ���������؞��*z�[�s��[sT� ��eJ=�-�k[`��z��l
�N59u0����
''@�e5����͝-�0�Q���$$
"���]p���Ύ�t�W���K���5�T�ǫ\.�gZ�T
�@��@�
4-�ӓ��f�=�g:S�r�̳�~�hv�F�A0�E�M*|Ӗm��[F�޲�Lɉqt6+�����C���`@7*R��Qڜ���t�����P�(gn 0��t$B�Fa$}�?F�r�^;����x�eZ��Z�D��{5%j5$Y��-��t��@!7$ ���P�VԤ�ᄒ�'w>�)��.ļ=�4S�
*�a$$B߾e�& '�����QW ��SH��`���[n�P����`��V`p��s���s�#W���r+��W���89[���y�9�j7#w�N��bCay�#��YON�%s������v��0�h�2�RIvJ���q;,xK��m����ՍU'�gB̹F�`��"�wZHEt�iXr�O v@�H�ڮ������`�ՙf!�:Ů���E�?;�}�cUd�G1�$��vUor�M��̻-2�j1u��Gse�1�ݥ��pT Z n���^`�uY��� ���\U�h�EP���w<�p48��@`vP�"Ѱ�Kh��H�[��E$)*��<�����7�L�twN�4 0g$�-N�Hm��0X�_�� ��u�n����JY���/I���(�i���N�) ��"��p��7��/�Ik�<x�?��@+AF�Zw���LӦո����
�8D�EuZ�<>*كHű}��+;��~��4]`�� �)���u��ĉX6!�5�N7n��l ��U���a�*@���1���Ao2��w�~R&�%='��B���~�&4�1�WT��Nͬ����h�����Ú����X0h�
�[-�NOcqn��)M@<�	SIlܰ�|E�;��p��1�����58z�(f�,�Vg�>� ?���Z��l��3�x-$"`h��(:0�ەN]�v%�n��[z��6����7!J���[=�( Ȝ �#j&���Ҟ$�E� ��SO�w�{���fn/My�;:/�& �սBS\�r����{�=���é=⚹&��c�$���N���;}'�C.%B�o+^���t/��A��$l��a���(��۶O>��9`-ך��B�V��̗��c�N�G��rӇw9
��(eU��f�]�TF1�C+N��]�P1ج�[�T>�i��g�{v[�+g���?e�����sw��h���4@��)Q��3������8��� Qh�Sݮl+��k��N�V��_������>ğg*��W��t�����/�|o�B�,NN@\��LZ�&2���J�\�h���B�[�R�, %�
�UB�r4�]�8-��D��yLI�l_�_�ڦF]Ț��?~���<1l�Ck����jb��E�]E����srP,�;��B�&S����+�?v����@�� ��{��n�	�����3���GS����e�,�N��4'q�/me�m��F�0-נV����������������I���w�]���/|�k��(H�Z�!�2:gju�mB$�-�,Wf��L���Z�����dں�T��<�#+�y��m��zU�o^.SqJ�BY�&�v���P�l�ڔ&��u�T\�rE9+++F�J�������B>��߃J��3'O�V-�PȡP(�T��3��K2�(�j��^����avn������߾c^�߃ѡ,���/�9�����-R�֭�},����G��q��Y���C��o���r�]��*ދ����������3|�{��HFE��� H�qevN�"��t�#H�È����������Z�]��+�M��h_�je�&
�y]�Eԣ|��{�L�R�l����@LcѧW�ۋ��'�y�
Hxn�sjJ��ƀ@�Y_{p-sM�`i���>qo8w0�?	�N��2$0=5���ũ�'p��a�	LS����	�mJ�ͅ�������<���
 ��v��O=�M�����>�ٯ�G΢�4�H� �����V����`71%'��)]��)촑��N�)���W;�Z�_��%:�� |҉5Ei�hT#�ɡY�u']��΄���3�+`Иuy5�`��I#$�����9&:'���Öh*|�:_�rB�W�E�/L/��U]���ID�Bս���3�-���=�h�,A�Y��^�K-}1��=�ݴ)�X���ν���m�S�VQ�vyG����HOp��DǸn�6�� ��Y��@ )�e�dG<�Bqԋ�Y�[$bRk5�����z�R���P�j�FU�nQ,��3[�
��q/ds�gP���7���^<����_�P_����r�QV�����k_��x�Ο;�V�"`��"5(e�����~��~K�G��7nƮ�L❿���g?�YT�5\:s^����	��DR�:,��L�����c���    IDAT�Ѵ	`:�'Sͦ�ZKs�R������i ���
I3 �T�=�M�K�Ȧ8�{U3��ھ۷���s�Ns�ʪ�t��_���/* ��m[��Wރl&�i��7ބ��Mh���/Ǉ�������}�,W126�u6�n��C	�NLN⦛o�̚Q,���կ|b�p�u�����i�&W��a~~;w����gq������g�,㓓�����Z�ܹ���q�ʊ����/�}�cHeG05��vKK�h�y�Gh��H��
�|�i���6��u�7s�J7��YQ{�G�(vv�ӱ�їz׎�)��nU��Yg��K�_�{��t �˟n��	D�{���j�-��y>4U�P�`���&t�1+./�wu��a!�]`�'�X;�7�gN�C@&�"M@@8˧ ����w�
 �w�)0X��x���xny�N� � 3�S�%|���GΣ�Pm�hի֝WћT1�vj$��k��#r}bq��a��]�u:��v��v��u*�F:J �27v�3霊�z��u�/IH��h��L�<'#� �����e�+�)��*��� Gbz��^t�'s�xw�Go���Z�/�//�g���FSw�\]�3uŝ�܂�L�^�h8��mk;!mo
uJ�ï���8g1@���9�{ϞՉ�)D�;�K�670��v��][����è�͙��@�H��nµ�azz��j�%4��S&"�:;��;`P��h5i����A�� ��HT-W0�c�9�[6nF&�����K5;~{o�'N�ĕ+�(���O��_���S'����(�,����p��
o������x�/�S�s��l�c���}������~��/`��e<��cX�a���:�$��T'�,۪֬0���L��P�T��34p ����iQl2Y��ڨ�K=[؞ق�(b˓h�zI
��A�l��;g���o��7����^~�nۏK1ig�J�/_ƙsg�|D�Sw�y'^��{04TФ�Uw�~ՙ�'y_L�Ƶ���!T�U�ص�8)�v��E�.�b��)Y��$^��[��f�q�:������ȸ�SN_FGG�c�N?Z��߿Q���Sg�X*�[n�k_�Z���{�t�C�_x�K�o��?�N��}��X.7PZ��y*�rN�"9:���(��݈JfTM	�y�Q�ݧ���۝�}B}Md �8�������%�Vg�,�M���+N�����V�	��q��L�p|ˡQ/B��> "����z����I�z#o*`��DSF1c���5��`]8��C6�E B:�p&��~��3x�V`�� ���Z^�]����..��!@�A'�����ғ'����%�Ѝ�h�D�ms�BY~[�ԋ�`�0�]-KȜ�QE.�ǆ0R$��#R�DHEF+b�R�`��":]�U+5��jXZ���$ ɠ�&U��f�铸�&2�����@)�E*��}$������&���*��[���8��\�\�F/������QlT��B�
!���D�ݐހ�2?њ�b%7 �2��v�n����YD\E��T�Ú���Ю��\�HKb:�&@݄�ר-P��n`��4��ߏ��<�t+�&�-~G����.֌��n�&��W����*p���gQ.�T�nؼ333�ŉ'l� 2Ԝ$*�P,k�e�\�|���p�
����_�ʿ��?�	|�K_A2�h��Clڸ��X�vF��D��ELLL���x�ч�o������^�'�x"nwb���[�ȇ�s�/*�nie�T7�|+r��v���cO=���2�oۃt����ϣ]���6ĴD��ˌ�y�S*��4)a4�G�&w�U̪v�V��	��Z�01�����ċ_��ݰ/{ѭ�z�;w1����.����hǎس{��u���F��v�}*�����{�Lp��lن�(�I�/.
�q��m* E���P!�l.�s����)L.��}iicccX�n�l��@�2�rY����_Pw��=x��_��޶�������Cx��� ju`��۰�\���
8�lMR�I�#cH��A��Z����b���Ӱl��
|��_��6�)�K�w?���*��w���uqy#���\p]Q:�=�3 X��؄TSM�K؄T�IW�BR��ǽ�G���X�}���V&"���Fp�U�����3�G!��1~�?�[v�*W�OŃ$�`���t+0  �tk;x���
p�T*��袎 K���W�ĉ���G�gD�b��ė��&K��t�! `j1�u$�ˠ8��l���p��`�q����2��*�D[ $�sQ�VU,���A��Œ&��4���[�bq����R�f�f���@z� �����A-q;A:��Dq�+�"�xM��M|������u�"��xz#W��u=�Q���	j��\x��F��B]����=\��*�-r�9�`���9�ӯ=�vľ Sqe.\|ߐ�9�l�lF��Ң��6Ϭá}O�~e�tL�V	u8ܳ6��66���K_|+^���156���<nؾ�������x��i:z��Ӹ��p��9T�%<uc�6oވ��9�8qJ�N.Tj����n߃V� �f��=%�B1�L�Ȥ9���"v���p��Y���P.-�҅��� mߵ�����c�Qם�݉}�k�z^��o�n����cO>�|�[�n�x���I�dsE,כVN�FR�T���ZN���Z�V�z=4n/�L�$RtX�iw��P1���,nٳ	?�w��^��o�{��/��Z���:�C�#�
���Z�ې�]wޞ������͢8<���r����t���� $�u�s0Jˋ�ˡ-
>8i�{/�+h�x��0~��o� ��6����(��D���2���p�=���?��i�>y�_���O�� �k��|����
�� M��Dɡ�M��_�{W}�!�ܾH����*н��w��3�9�yA��ߨ;rnO����> ��~=Y��	�6�~州�ev߲G+��P���ξ؃�.��o�.����5�%��4u.���ؽmN�8��K@��6~�����"�/ �l�{ny6�}>��<X�� ��e|�w�
9u*�_)�T�K��Xk�r���8��y�DA D�
>��&�I��U��"�6���Na2F.�`�D�����H�J�&�q�8
�F�X36,3��|��/.�T�a�T����pqvNm;�D���U�T�1�\Ǚ(��&�,�U�vH#\P�=ҩ)�>P;�D�^����N��}�
�Ɵ =@¿zJ��j�t���r ��X���X�&n�&�~��IPRP�nW�������xeV�f|uw�KQmb��*��A���]X%L{��5D�ٲnG�~��9i���&!r�j�UCt�u�~�5/ŋ���4�a����|�I|��_hX�a��iB��r�b�J��\;
��_v�K�*������Aߏ.Z��M%�JyYZ���q%�+!�R����{^�b.����,��ݿ<���}��(��ظ~��܃7�ؿ�j?���ߍ���c�엿�M;�"[ǁG�!E�cq�fV;��M
��\Ie� ���]}<==O�]ݤ _.���H##nڽ?����/��[>Ǿ���1׏a��P��vddȨI�*�FFu�MO�����5��-_O��/�H�B�bn3�!O��)�ә�����s��&j������_�˷� ���Ii[��G��TF�m�(����Q-����j���Sң�ݸ�N
����39s�ȉ�!�л�G9���{-�4�p�H��$W�I�kB�����G�t���E��[7�U����@��l�%����M����:F�TWƦ3����)Kt9
2�ѨZ�Y�>ַ|} �iں1< 9y��\F!"B�����mj�P�K^4�`}�>����� ��[�m\��ǏǳK M�h$R�����__}�����"�i[��V���2/A�0��1'�[J6��Ȅ��8���'�A�d{�m��X7�ڮ"���$;�^H�`�}��\��0�2.�-����x��'p��9�[y��A�f�O�b��B��&�}�\2�f�*��,4:�{g��
�3�I�@��!�������(�/��f�M�����=��v��N�������M�$�b�@ ����,T΍����5z��[v�I�ݦ�9n��0F�V���\ӷ�Ï&�r�y�Hq}�6��F�m�ǁ'G�0�(�E:Y8b"@�
e����غao���=/�#��Ϭ}6 9x8>r�>,���(n��F��,!�I!��aiiA4�Gy���
4r�.��$צ��E��d�h"��v�
e�fQ� "��6Q,�%�&���1�Zo����7߈<5'�.��+�%�ğ��=���6��wݍ�k�arr�6����7;~��~|������[p����7mrGp�q��%� 1j�G�
�9Qpv��"�搓SJz�\:B*lcl,�W��V���/�q׷|���W�s��t����T��R�6Q�ΉH�R�q���)��lLLL�o���|$���uAbe�O�J�e�-�	��a��y�c�#?�#xӛ�$`Ó�V�t=���8MmN��I���C��/}�+����86���bv����U�9r�N�b��<y�{�(�t�"[@���I��� ��S�\e�I���V���� �ՀCA��K�����~,�z?�� �4&Ҥ����N4ϐ���� ������,	�g�9 �c�v�;yWf/	��-��[_���nʳH�5�s�݃���||�k��x���O8�$t&�W��F9,6���_���.��N��̠So��I�]�ŷ]IY;�Hu*(��g�86L0Q �Lgp��-�i�VdC�|.b���Ta�m6P����i��QG/�R
���)Lͬ�Ć�7#��u����w�/7��D7���|���o�?%�ʌ��H�Ѥ�7�
=7 ݠ�ܸ� �|�\^btN]��P ��$r��v�,�i�Kx�ߚL�VK� N�l�Fs95�-U�珻J�fAL��0�E�QG�̓�~b�19��ҁF�L
��
rCè�+��3:�L��R
�µ)f'ЪkZ�N)�
��(�B�E;����h�k�mN�Җ�U6H`zdG�=%ke�4��;n3��|:��^|�M��}^|�M�>5���ؓ���Ǐ�����n�X��͛Ѡ"k��5�X�����Q�U%�C�bu���^�����G^��Y�4���vyaA��E��~�2��z'v�ڮα&���[r���W��cGOa��=)c˦��R�^t獉��_~+>z�,��/�܁��'��<�TM�c��O��VW/U���Z*��e��a��`�v���Yw���h�ҩ0+s�b6�T����!�r����?���ƿ�s��/}5>u�&&�`iiI9�֭��¼�btdH�J�Z��w��]�����^�2�bp��7�Z:`nذ^ �u�{*�:>��Oi��oߊ�n���wΞ=��kע\i�Z椅����0&��q�Z~�cÁC�%&_�n�������AG��g�⎻�ƿ�����&֣��an�����uq����e@I������o�[)�!��~( �oa�]�\��
}G�z�[�ZB��-���u��a���Ż�=Ǉ�����U��3�p>�P�UM?(�oK_B`��M!��F��m�V,]Y��cG�Sȅm��߈�� �Z�P���7��������� �|���?{�|j_�R��s�L�h �ɹ2>��'���s(��hǑ$G}��A(����]C�[��P���Z�=���w��mk�._�Ƀ����ʑ��R����ۙ�� :�sc4�Eh�;�֘���iB�/��{�yJ<}�0>�/��|��uX('�P.�7p��<�ȣC�.e2�����ìB&H"Ȥ%N��7��:�В���M"��>�ĶւnQ^ JעT��Dae⩳a�֖�d���.���W�G�'�)BH� EŖ�N?��[���B82�U�HD.1]y(�6���7� ��O{�Lqu��]!�о�j]b��$���NA���\�/���B�l*-q2�6�ݪ#vp����7��n|�����뗾�H$�|��@�ڵS*9a��b���}�� I��ӧ�bjj��7��`�R����ַalb\���ɟH����{v_���?��O�Z�`ff�J���_���0���a��5�����|�
6�ۀ�O��ڵ:�v�مu6���S�]\�?�1̖jHOa�ݸ<WB����������	tk-��$SÛ-N|��\�8>i��`h&�j"��Hs�*6�Ý�������b���s���'�'N��¢��&qr4�uj*l��
��|!�I�k�����ڵKT,���7�ᇿ�?��?�u������o�W����_�Q������W�:���=�>�G��1���u<�y�k�K��KΌ��V���I|��GqhgϞE"Hk�B��cܨ��/^�z\���3���p�翊�'�#Ne&��4 �$r6Ho�뵧�hX�L��U��Q+^e ����J��kn��dx7���} r�������[<�x]�	G�K,�ݜ�D�������><x�?]! QcE�=�_W�uS�o 9s�� 5?��7��6��*^y� �pPGV�� ��]��߽ W��}���� �j��x� �:v	�ݦ,��?|ؖ���H'H'��8�n܀�~�^|�-;Q_<�O���(/ �HbblBZq��Z�|j�,�ȿ����;�u�_`��0�m�߄��;0�y�ƣ����0<�	�V�F
M����Y,�;��c��9#�S�Iǲ�:N�k�T��6��I*s���8j�����|']^�l�x(�#ف�ܒ�:��'G�K�٨)T� eH���d���n8�)F�p��q��+Ѥ�T](�hZ��-�����Ӹ�0�Q)��O�a�R�K�N(���(�Z�Ŭbb�۱hf'=C�Mi4�x�"P�H|��Ď�#�!��
v�X����ރ�߲񯽿~���Q*�n8'!;vlC�V���� ���?�au�I/��Y���������O��q�J	��Il[;���SW��{������߈��:���˿��� �'��RZ����;X31��K���$Ǧ�e����g?���"�����Sزe֭[��o�	�t��!D�؟G�^Dqj^�?���+x�}ظc�'�Q�Uu.�y�� �|�� )�afzTK�Nif#-��eZ$'�Sױu˔ ����ǎ�������,5S+e�.����k}����J��L&�x�O��~G*�KNM���w���oWP���cx������д�O?���?���Y��}������{��~|�c �ՌN����׿��x�O�U�x6H��	'&�w_�C�������Ew+�s���o��=�ȁ��J���W����h)T�M�;-	�I3�9�C>�ZJ:)���� �ht��G���x�J�bޯ��
ݟ�`�m��v\��q͟�Z|;�kO����]� sG�Y�p�~������~�.�+r����?� a�Ky�$ �	C�������݈tk��^�j�d%0ةo�
.�o�*>�y�ǎ��//̡Ro��%������Nϡ�ɠ�H"�%(�ݖhGt��k�e�&֎Fس6����a�T
��S��?���F��U�5٦�\�.;��CW|}�\���H��t䪓
��U��R=�n�������;������O"��@nx./�8u���$�,��h��dS>t�va@�E[v�z@STF��"NEh1�O'0��_�J��a�me�����@�7K���e�p(�=)VS�]�����[7�M95Z��&Tnjb®)]���a��&�	�0���֐���%NZ<g���"% B�Ddt�Va��;�4%��uZ��H��Vĸ�N=��:��r˺�}3���씊�b:���c�����    IDAT��w���oMzj��x߁}h7k��Q���{^*�$1jX,s2�k��k8u������~?�C�M<����~��q��Ylڴ	O?�ȳ��w���?�l]7���SO�������h�j��?�l:�Ж��J�(U������x���B�I �����ƍ�뺝�7kx���12<�O��<����l���^̕[8p�4�LO�Ѭ�Sv�G�G�ft���q��}@6��ﮤ�w���|��t��$'e2�hR,��g�F���m�O�~�|�9�?�8q�t/�ZYy�lV��E'���D������ˋK������O}��_�{��^itΞ��8v�������}A�n�޽������C���p�2weoy뛥�V�ѨI#º�駟ƞ=��G�O����n��6�ݮ�;p�-7j?����s�.���~�?uW����.h�L0�*\���P;�k�
�O{�ѷr=���+���d��\�_�������ȷ�dI�՗���e�PV3���ĽNS��M�G�
��L��Ԇ��C�v�l|��B�|�_[��=
���9�(��H6��yӏ����i������w@�Q�k?�3�3�wUVŲ�{�el�fLI(IHr�KH�q	!��C35��F5L�Řf0��Ȗ�,Y�յ���ٙ���2&���Mr}�t�[�;�����|OK`�g��̷����������vF�矾k6l���y�w;�y<�r=dMg bc7��5 �K&|�"nu�jpԌ�ϯ�)5~��X��J�c�5|(�S�i9#�	uthv��P4�[G;�d�v�d6�R���IÜ.�K%8Ag��=q~����Z�}���k���FދXZ��?�b�Ihה��d�u�n(}	�
h�*`�TPجE!����v�Q4��M\�\0RI~>��:�'��Ii\����!����K�P<*<��l�= �*�{��!��x�@�{���ڰhxdOI�
B<L'�)�+¡xZbP�	G^AC	i�s�]�u�(G8b��+$	2�s���N�K�d<�Xk;�C�@�Y"S�$d����,P^���7^�c���kGc�x����f)Y$�g�y�&|�kg"�J��ъ�|� �A��_>�t��K�3{ۮ=���OǮ]�8���e�H�7odZ�7of�'��կ��{���kot�7\{�t�57��>�����e3H����a%�׼��kX��:�!s�C�$�����o���v��^���{x��U��>�� -t�ĳ�f��5��������\VZ��c�c�{�в��c催i<Kj�y[����O!n��7�ݦ� ���2L�8w^��������f�L�t�y$��%���ͲF2�����0��� �%ǅ�a�7�-��n�Z�))����g@r�=�b�֭�R��.�cƎ�-�܂�^|a
/��:�:H����|�M�Ivs	��ӈ���2�[�q�\'MF4Z�=#�G�F���uǡ�*����xku=,͇�d��-z���ȑV}@��E����Š�b�ܟ� �;�bZ���|8|
���g�����?:F����%bD� ��'1�}�Q�x�)|E#����=|��:��¯��zJ5w:��,+	�L��v��7$�t�[_9	u��#2p�Y5w���O��<���
�<��37x܇d�6�=�^ĳ9 �KE�%�7�`MC+rR9K�E��qYA��B��(�QR��p�8n�8$��GK�Z�����"�_���(~nK'	K��I�8>�ŭ"cdy&��Mɲ�v�4|�����-��/���$RY�w���f-�����i�^(�*�m/�zs��K؈g,�5?Kz�B�aB�7�;��c ֽE�`��MF��K�hh"���f�I�`A)䐍����@W�H�����\
To6�2u�KAD9�����}���X��!����De��_�$R���v��O���0Bғ���o���v��b
��4�Y�E����-�g�n�'Tu�,~�̚>��
TZO�+z{짧�xؾ��[��'�cǶx<~ds&�֎DWw/K��l]��+.�9g-���׍oo��
m�K;��,۶�̳Ng�?���}U�����U8��8�����N�睻`�X�n�ο������6�g�{��v�Ϝ!M�;L���3�]y�����{�V���n��կP[[�g�z���߉��_�=���=��_z�ը��Ĵ)��#d-�����@����b����ӿ���8�Y�	#Є�&�v�Jg96������Hcݪл��[p3CV`�����\gĀ8)�
�yæ��!����c���/ָi�nALR���{�\�ȣ/CI$���J#PJ]$�hFl�O~B`/�H����w0u�4���k6���@rʔ)��?����Q�y��eQ�~����x��7��?!���������k_�1���q%�I� n�� ����������*h�}��&S{��O	V~�/��J��;?�3�ⶩ�ؙS ':���������[��,���;x�g02�����@���+~���z�ĳ��RLۣ��墴�9����@�{��Z)"u�8�;����+9
�bi��)��x2�~/��E<GkK3t�w!�o~�xQ7���.rX8�np�:$�ăO�yX�����p����z����X��@��#')�4l��a=V�݆�L���t�w7��+�������r���/��IS�+�ｄ�[⡎�Cd�N6TdI^${@�˾@�eQ��#%P57k�3Fv�D_o:�[��]uA��B#	ӈ�_�~dEC"�ð1�q�����܁˯�ޒ�(�K��+������,�������@�mf Rp&nj�.�r1��P�;��:��1����6R��I��y�0|HF��hm���e����B�!/ipi�q��ׇ|��{g������n�o�x u�*"�C#r��K�t�;Fބ�O�Ol�����=�\�2�J��+a�����+p�2���0jh?��`�&@wQ���ui@��jUᓚ�s��L�^j�O9�����-[�lٟ�sW3�G�C���d�7MD|l�w�~�:�Nھk���if8�h��5��QQY��4`��|������u�8R3f4f@�.���Zݚ�נ�e��i��d���|�)x�e�CO<%�|j9.��B,:�N*:Lh.�jbо�o�;n�~|�O�c�=�#d�氃���D�Hi	�%ex�����o����7���BIY)#�_��y_���n�����CϮ@Cc�P9�S��<�N&I�t� f����`՛+��A�za�(�������T�I~��-�ƣɐ%����������_|�544J�J�S�<��ő�$yW;-�u#�9�l�y�@+�^���1������n��z;V�X��3��B��_��6N(#�:���S5��۶5 �La����j�z��h�d)�I'3o8�k���'�Z3K�L��Gík��V1�B}@��ڲ�����niD[R C��l|P��z2͑�H���S�����~>�C2&g�h#�d��a�H0�x00��e�f�"�P�_<�_A��� I�@���6�������981���4 �^>������X�H�"�[�xu7o~$��h�/��f���'��ç�e���p�������3���+�9]�A �9=�o�^����
�V��~�7�U�a�%(H:��T��Z�EF��y|�~�ԍ	���c�\��d.+�냠4'*Ȓd�*�˃��̪�_ J�q�����dϾ��}o#�;[�{PԱ�7@%�^]�ac6�O�^���x������/"T9})�]z�6�u%�j~�s�����b2ɤ�:|%��	,I��8��h��+������W]��p:a)�uIZ�i�?.[��~�5#K��܇@0��&U�`��f�p�	�p���B�τ.Q�<�kl2g9�n'0�i
#��d�sG�6u���=��/���xJY-��I�B�R���q58�c0m�0TDܰ2i�!�uF��S{B��6�:$�n�/*��yD"o�����翼ɜ}���&y'�F�'���7�E��[��|6��罽}رs7f�>G,\�ݻwc���� �∅�����k�5���o���ˠ{=܀����Ǹ`ѱ̀xy���;������{p�����'�(��4U�����`��:�x�	x��?�iw�����d_��'��DPZ�3Ͻ��^_��?�1��ƏCuU �1v�8̞�����b��v<��j�Jk�xB����)S6d������9F�QCj1�fV��6:v�(����\��4���i#�F;�bpȓw]�����;ɨ�k�Lg��z���5jj����B���$��x��w9ъ���W\���\}��l^B�߶��6W\q�.]�1�tވ��l���(-+��D*�_\r)^x�%�w�o ^t�E�]7�����>���@ee5��0��E �c�bs�l��1�}����zГ�A��(�ur���p�^�]! "=X�b,�biV�SGPS�S��)�:�K�ǀ��Y(N�� ���B�S�f8�q<����gfx��t�}��/���;~����,FH�2l�� #4�����1���M]���!�[c��B ҉4�[���? @D�AU2 ����
�+0@���|��
��\/ۂa�L{c��ڊU�ї�<P��(�iA�S�e����|�x���=��S��������^2d�� ��y�Ce��>j2�
���7݇>xA��v�<��y�:r�0�).��ס]�,8v	B��p����_6�AG����b݆]W� 2js� � Rk����@i92��jl&�J��9'B�z�>�4��K�=l�L
2����kЇ����ۇ�zS�y����z v���7�l�u�w��p�R�rIL�$;�o7��k��0ƒ�\S�q~IjH���`>�9K¯�y�<�&D�(�l>-�)�w�_��=cUI�ٓv���!=���+|}kL�"��KRsF���>��eI��B6��b��Jx�w�ᘹ#�w��@�S�\HR���v�Q>㬳`L�}Y�~-��/\����mJ�A-���s�z�)f%R�4ZZ����;ĩ�}	�q񥯜�'�= ���+���5��n�s�פ9�s���Ko�5ܽw���5���� �f?�(��X��T���jX��{xo�j�u�<��BEy�>�%*�8�����}⽷?Į�.�����E^V��܊h��yIFO.���B�<����<rֽ��I�Œ<	*��?x ���B�
�q���,�1�n���ҿ�wv��%����z�BEoO�=;�jk9�+��C8����	���7�{�=, �	�\|��h����7�Ma��Y���p�UWc��u�����zn/$����{������o����0{�y�I�.J�6)#�Gy�T�a�1
��J�����ؾm�{֭�.�5����_
A��Q �i� PZ�4��h�$�\nVUJ���I�vB�0U��'bS�1a<�`���"CJL�i���d6p��t�|
hY�@�E�B��Y�P
�n8:�OzH����֢��J�t��
��+Wds�*�M�l���ql>'��@p�'BA	�Xa�PSU�ޫ���̾������X<��>D�2����7}v�{~c�����V`�����m�Q��+��ƍ°
�]*��}}��؅�;�1 I��LO�H�\_/�^�с<��Y�Ɔw���-kt��,M�2Ñ�\�(JkF`؈):f��}�u�lM;7Ã$4d�ذ�l
:��)nlol��98��/�[�>)�-T�XZC�P�cOlՑ�РE_�d�^ލV=�E�%���AsEA���[���%p�)�a\M��Z�P�6u��9�@c}�����������$ST<HM�2\���`=��q��9�����B���F��J|}�X��:t�ln�A�v�'���f���e�����u��aRYPzf�.q�O�=�p����6\�H����ݍ�2/�|�n�zH9t���M����u���$��]�2e��|���eƐ�t��W\7l�Uѝ"EX(	�x⏿��VJ���B$1��\2�{z��ٍ%�/FKSƌ��][�l�ĉ��A�\T@ig�(n��v�AX��62I�u3~�t�c�N���a��J�.�E����`ٲe8f���}��z������w��~����7�l��=�GCG[;_�Ke�6�¿���X��&����U���a_ ��$QѼ�O����+/���1�����U|��`�эH8
?��r��q��>�/�-o-�w#�H�'��%	�bb�(!�Jb@�B�� �m�s'������P}}��� �N"O�Z���H&:t(��T�>���e(����{[p�׾�1c��֛oFgw7n\z=��	���������?�9.��̀,^rK�^y�\y�娩��7���/��2^~����e03f�(� i���e��`Ԉ�7n{GH����{����֡����_I5��`i(1{ȑ�S<w���ʐ!���2'@���:yȻ�a4�<�bR� )ʘHL�8�!�`PP?��M1�����?E��@�%Q��uɋF�E�DE��`��A�
����]�>aM^�1�;?i^���X!��@(����Cj��% BW�+��٧�%ĜoGH��`�̿�3���+t����jo���2���ev76q/��a	���:�~Wz�22T�Ar Ӏ���6=%����oi��'ź���O�p�a���B�u��
�=�'Lǐa�x�U6�(6�����6l���_S���5(�5̜{^x�m��x7�@�AwB��}������}9}K#�|�E�Wh 5��.UA!G��l�*ø�g��o>J��)C�;)�זI;�LA���|� �^	�_�+����C�zKaB�`������e���+!�$&��w[�ĵ�܇��� I��$�2Ѓ~L;3&���'��UH�Z;z�VG��Vԋn�yw��`g�q�	�����@���%>�)'�.�=�:��y��E>k od��X46.��o��Z��>�ڑji#�5���t��_��4^{�!L�>X��h��Ȼ�4���96Yϝw֭[��@�)Z4M�����u:Y��1R���[n�ʷ�f�tWo��v~��Ŧ1i�$|��C���
b?~���qʱ��sr������w���*5��7K����Ǘ?����I?�V)���`8��k�b���4b�fH-<~C�����! 2kn���$���焿l������Pu%6n�"i�I���+�`�Qu�gV>��z�;Y�'�Y��d�&���f;�w�Ղ���it�n�0<p���{�~�V�����92���!�1�����Ț)f@�xNiW�d|��j\x��;w.n��Vt�tc���|~��׳���:,{�i���~[��|b�<�L�����H��]q�fKk�����#n��v�i]s�5���t��$�εA�5˟|�1�1c�M��瞚����~����z<.��E:�D�\@�6��lx5xKK88���  �:O�9��|��	)�����n�t��P�ý����8ۢ���)���wC�����ޢ9����|�N����A��YH�� $������'�#���Ŋ1*b��v���D~ӣ�9^�î�����$�(p�9��Æ��?���{�W$3��	�f���W�|^���yhV`��u|���
�ok}���C((ߩ��+��F}k�I.=�\&a$��%�h�0����$���@	������˭��P�^ ��Q�y����s��o�L�~܀�a��(�9BA$MY��^��z��%0)��8�ڙD2c��'#&}�79�.d.���    IDAT�G������0M�6)�wδ�8���1fXFTJ�u%!��-��òǟ��SN:��/�w�D���Ql�ۅ��?�7�]��P��8i\�i!�p�Qu����,���]ۀ�|�i���x�~���[����|]���s�c^�O�K��acruPr�;S(�J<a�u���e�� �D���ҋw�ǟy	+�l���`)��g��K,�
��f|��c��@��A͍�aIy�P�QnD�����*���c���#�M[>f.]�����ZM>�N�l�c>��T~�<\Yn�Fb��o��.���^��عu���e��뮻�}�R�ֽ���j�z�ꫯ��h�#���<K���Ĝi��_\q-�Ej���ܐ-�=�'@I�M�8���!�5�x��x�Q���G,`�uyI	w��Ci���0����p�5w�wO�	,GوZ��ol���{PVY����!{V��B�0�[;�[�Ԭ�"�HBvbj9���y@��nj���f0�[���fO���۸���{{�a���>��w����$ݛ>u*�j�кozc݈D�z�{����~�V���Tj̸�hmه�3�sW'����Gɥ�UUU����/��������O����3f��sF�Iᮺ�
<<���t.2ʿ�����\bH�ɗB�gӖz,��V��3(����1Sм��}	��t�	]qC�x��C�PY6�^�<Ŵ+�ӋigT�)��0�ƃ�l {9|��N��ɡ�p��XU�ՠ�!y���Z�a��>�.@u
���4���d�Q��f�(Rl�w�)�A2.A,P��(<��G�Euq%�	�,�s B�ՁOd�рk��9����;���=��7O;� ��u�����W��a�����0�/�~ap��8�@Ց��ص?��VmŞ��M�KG�?�ѻ�TN9|�^<��M���5��
��tڎ~䄌Pi-F���!��?��̾Fѵ��X�N�'��bs��S}A{�7���O�OϿ%2
�B���]�}HTpH	0.����	��~�+*�-(܇�7�p!�l������?>����=xt7K=�n��?>���{��§L���~�L�p&����b�а���7�v7�x-�z
5��T��5|�ą���iѐ���O��
j�q���?$f���°� Zvn���BMH�[XN� %G}UDjơ��ê���1�RC��ӇF���4��z)��d��2rN,�Г���\�{)N����S�-��P9�stE�������C��2���E&��`�G�?�>�ԔMe�{�4c�揹)�����TlG;��{�G ��)���s�=����5|����؈���Ǿf1��	28��/�{��k�>u�W_�T�pݵ<,?��r�)����x����HY)^x�%��Aj�cɉ'�ԫ,R�iP�}��Ӊ�X�uu!i�ўʣ9$�
�}'k�L��ш�CG�2Z��H���LZ�����!�Xt\�P(�˓.G&�-��
Y��,��<���\9wTZF�㙉���-t����i/��KBp�����P^E[gb����߶o?V�X����\9	RԤ^^Y�灮��/����Cq���.��ͨ���4��B���lb�ƌ�K/���.��Mg��{�]X��#�1
��D�>��պ�?����Kq�\��Ih�I �&&�v�	|S� ><�L�Ql6�E��@O�'�<5"��{�d|�3U�x*8���S���|sb!�=$�T�$�:7�A�^�w;>��0�8��*����Rlt��@����t/�c��B�}������_㤂�g]�x�����D��^�7F���l���V_;�h=o*#�\��ك��w�����?�>�+9���-V�aw���!W�Y�eM]�x������Y��&t.d#��+�������/����B�u��VCe%�9���Ĩ�31t���YN��.\_�Za���-lZ��m͈�G�ɦ�f9w�b(�r\x�-��x��-{��Tq_G
u�P�JY-�e�܃B3�"ِ�$��Ń�݂�5�p���JK���ڋw?\��/���9DKJpĬ�8z~N�;\�֑BU1��#���%�}t9V����Z(@6�q�)G�眎d���R����pߣ/ �JX�n]��lNΛ�	M6!�z���a�W����UaiN��_��&��(�����,x�F��W��?��:t�����4�:Y�4��P%$�
4�?��i��O���{m1r�Bf�b�q�6��~tm9�x��3�R���(���Y�ʘ%{IH���gBFc�	D�,����&���؏>���8!�����=O�߹ML;�?�_�mq��7b�˯��7u���ji�Vq�Y_��߁�u3>�9˯�7�p=���K8��/�˻ݔ��������n�ko���fb��i��-d�#A����kؼ�-]]0( �����"E �녝���z��5�e�����@��6
�z(ԁ5��
9ixT�,,�.X�~��,$��T$ه� ��Esf�ʦ��ƭi�C=-MMM<@�{{0r�0~���h�ꆑ�A�j�flٴ�<�Z�[�\��	P�&F�:g�+bdr,�Rd9�<�Xo�y^?�Ra6��b�I���h=���r����R�֛+���	�QZ^��a�IA~m]�ࢋћ0 i̚����/��~0rs� �@&3*����n[α�o�$X�#�D��X�QL�"�Qd��`����  M�nA��=!���@zށ�"(`Ef@�9䢷�7;���|&$�"�]�T"�	DIdw���~x�X>HFs~/E����<�>�V���)!L�ܐ4��)��K/7 �"ΈJ1e��	&��Z�߲�S��|�/Y�#�!��&p���3�?�6����
�<��S?����
�n�+(�� �%)H�7����	k���7Kڵ����9W����:d��aDU�S}2�� ���1u���:��o���E��	��v�7mA[���:4ME�̣v���1w��OX�Ѕd!�>SG*�Cs{i��B4bl8J�= �4
���_�~T�X<o*�s�I���Ȥ㰅������^��^yݩ<$��,�eJ�M���r4&��E2�@��*i[J�gW~��z�,�S\���q��q��?�^�q�~�֗?�/�O����Y������n2�
e3���{�1�1^Iڵ�S����&}�����$�Q	⦫/@y@�^�0*�^\�W����a* �Br3;��B�[�Q4�eQ��W�í�t�6ǅ;�H(�r9�=2����z,�2�w��z��OB�5�S��u��#�\<�$4����m�>� >@��7^)�j˶z<��,�9q��8�̯2�����;����x镗��?������c׮Y���'�t*���C����ذnoSB��_:���t*��y���G���^��u�0r�h������fx���[�v�D� !��B�T"e{��@!>/�``	��%M�"o ��䋦g��P�1N!���@)K4[��@2�M�H�(U�ݯ��q�!���\`dӜG�9E���{�N4�ڎ�Pcǌ���a��Mm�tQ��o����Vғ�3T��p<9�W��,���Ws�����J���_i$� �p<�=ɯ��P��9�|'��i�I���g��]X�n*k����
�ը��E��F~lo
�=�����b�a��ع�6y=T7��=B�w�dR��PZ�.ŭ�2k[�u�AބM�ŝ' x 'y�bw�I�D�Q��_����*�OҤ(8	S�	G:��s�0�B �h
/�*���=��'T9ŉ����r�"�T9V�&/팘�_  ������\�|��YwC�x �)TÅ�@1Oш�9Y�đ���f�߲	!���ř'� �gS�G ����
��+pH���`7������*b}q������z�5;�P�������x��׆q�Q���C���"��/U#����A��>3}���k��="�߆TO��lA{�N�`I��Ջ�O=Ͽ�O��WiFgR��3�> y �A% �ZZ	����|<��r?~z�8��)�
&l+��B_"�����~�MԎ�S�p{�l��n���|�����epۤh�������C������}8~�D,��b��~L�F�;߬�^,�yI�vt+o�#S���;�$)�+��s�jSg�QQ.�=�?��G`�J�~}�E�
�n���Y�S���Hj%��ֱ"s�E�CQ��f�A�t�\��/Cd�0��I%Oi/�#�Q�<L�/�7Nvؒ��fA�ؔ�D� �O(,hA�M��dÇG:��5�����&@�񴣞��8��v��qTVU����Y�h�����������ܚ¯C��EK��G.���K���C�KC{Y����V�[����b̘q,٢�%�S]]�_^vZ;;a�.�"����O%0����&9���Y�M��J�ȷ���X/<4�$�$4E���#K(�v�P*2�^��#*�t�l�.�N��K�<2dE����Z�ۻ��"�%YS����h��!pGiS�M�>~zzz����k��|��H�<�Z/|>����<R'�#������8dH5��'N��8a:��;٫(	�N?O��m�������;�[����2�,9��oEӞ�P7�@�ʳt w ˥�= @8Y� ��`N C �3�#D)X�Y�Av����H�"��[X��sA�g�E�|w�0РD*��(�������7���x|��� ���+��썲��nG��t��B�ف� +�"�$�Ę��#'z�n�t�z<���G�I�%�Ek�$p !oU�7� $��A������1�A��`g��x�C�����.|��8�+0x��|���
,�*�n���T�~�q��&�}�1��)���.ł	�!c��O�ܣB23lHv��(��󎂷���u��P�)�5o���d�}KCfAR1c�h�3���.��.C^G_ރ����3Α��3�BTca#\R���%�Yz)��,�@��=��)�a�Ē:z��e���=�������p��ƋD*���-{����@�!��ȕ����n��˱���q����kaZ+B
�@Hb#{��5J��q-N�vw'ɫ�Myg�(J���((�.ܽ�T� dٛ[�Wߌ�^
C�:C�����F��CS
�Ki\}����I����]"-�P܅���j\���PT!�)�-��sӴ�M����ކ�����|!MUq�i��2�A�#���pQ��h`%ӱWsz'h���$2�n:�meGH��?�^?�l�YXSe��uC׉��בq��~�)S��`N^�Iz���ʷ���U쁠�ښڡ�0a�ְ�8�?�����!p8n�Ll����ب��(�9 g�^Yb�¦$
d�d������(�{�>�y�]lڡ��^U㡔v�u�D"�S'CmE����v!��#�L"�1�j�~�`p���@�&�Db�B�lߵ�?�����(����쁑��r%�QQT$��f�����xY���R���A��Ž6
��s=��`mѢ#�5"�{M�L�:	�ׯ�˞D*c ����4T��©a���h��e�V��&���)uX�~3b����pj�-����A�� ���T�b���#7!Y<�"�G&� (q�d�>A��?��&ψ��<�S�?���Lԥ!�e�b�p�<'$�s�|���HѶ�'1�N����
�9��ي"#A�1��eڐU7l� IV�Pj�� ��O�*�{t�|��XBH ����s&����8��@��=b��T��s�@��6lۺ� r���qĬ	@|��E�{@>S_���/�� �_�t�?{�m�!z��$�`��E���Ͼ���&�`5�zS��ꂧ����C�hb)�W�����K64A�U	�/�13b�g��,�#2�v��$�6����LR�n�Ԏ��@Y-n��Qt�%���s:�.t�N1g�:�;؞�B���H�cXD��n�U!�JI���4%2°�!�/���L�@����`��riO<-(�����^\��~	B���(peb8c�\\�_g ��7T���~����j�}��M�FքK���|� r�5Yp�FG�+�p��?D����h�����ŏ��	1%������;��j�O=p��HͽIɍ��$�^r�����e�܄~я���׆\00�*
��E&c���]�@WG;w�܉Y��g?�o."�a�Y Q��w��+�����4Й9�r�adr����ɏ�A�v��nݑ�8���h�/-a�!̌,�����~_�c~ɐ�����ю7�z���'L��/~8F���a��*N?W]}-�;{��H�L�5�77BH{8hp(}��Ԃă�3T�����֭��b@d�v��7L�T���hhU�:�<�G�� ��PDA�ԋ=��Bs�k2��~h*y/��8����`�u�BS�.�tv1=n<���F�h�� ����cť2 ͙G�RWL�����f�Q�ؑ�Cj��ܸ9���#D��\ҹ�A{��٘<y2w���g���x�wp�u7"����<��)<�2�(	E���%�.l�߁H�0����}Ȧ�Æ�i���+�"O���d���|��DgSܱ��m:�uAw�cJ�99��C@��fѽ���� �)3tbl	��Q��UބD�ny#ǌI���;񿂙Vb=��˓��@��㝡#E���fT� +��E�J1�E�9aJ�R5f�d����/
�N����sF�\���B,%�q�3�{*ʣ�9s&��v`�����DX�E ��ic��(���=u�!�l�g���
��y��>�gn�7���4��r'^u�-���V|��	��ш%����BP��i58rR9F�h���K��.X�K��#��sN9��Y�g���;ᆉ-?@��y3�<����o���������A	V�3M쎂�>'���DVɛ �޲jd
*���y� K�� 0�: ����E�-�o{��px�I�j�Y�v�,@����7;�[F�vK�[zq�7$��!!ً�f�ů~�}��	x�A<��Z�p�0�0�xCǖIs/	
i�sY����f�4��& ��������7
=�7_��ymL(q$X�9�עG��� ��*�GlI��/W�o.�UJҮ�1!$M-�8�Գ.
�z+$	���W/`�(�܊^]Y΃"��ٍQaG+��Z9�S� ,�����2F%����mH$�<(����2dd�5ݒ�GB1�X|��,�?�KK#Rt�*q���Q��:e��6�0�$�0m���ؼuV���Ǝ�������9����<�"�F._3f������(��L�����8ǨL��$�!E �I"��"�O+]?��D;�T��0"8�����r�5����&#Z�ǫ/?Q�Cw�؟����O ���$���M�]m���ɸ��дw/<���CO�o����:35�����ב�H�,� �F�$���j�m�F(���� �<A���!�����1k�,TTUp�ȴ�S��G�{�G�?�l�
��sXUQ�7 ��f�jɪy����R'�j�h/)̀��>�$�#Y-��sB���D�&���C���kҋ��N����`�a��<�&��y<@�(��9ي���29e�r@�����&�8�2(l�d B,a;�,$G#�G�>]��L^��i�0m��h#B��,#���l���b�K�
�sM�@��0B��1�2,G�X�` �ܴ����R������q�a��瓈�fL{H?�?s_��<��
�<�b���
45��X"�T��hQKҐn��q7�_���a0l��DC���ӆa����vt5����#�s#o��=��1�@ͬc�}����6=6�]����,��n0�!�}ı������)P��~�^Ӌ��ƿ    IDAT��#� �IL�ϋ@E�B��,��p�.B@51aHPڶ�C����qeaiKG�0M�j�J�:;��A<E%s
�GUiK{��R�����Ssc�� $� �ق��q�헱��헱rm+~v�m��ʐ�^'Y(�t.D��!7�E�e�����HҎ�>�WĨ�2i����!�20vX%n��'+Y>O#�%�˛���]rz
^di�~���v�9�G��JJY<�Ǜ0�L����bx4 5v
1s��p�C�Kd�xh<��Q�)�[�P��zyy9ܱX��>,8�p�L�yO�v2񸓲D�8ڻ{ ��t��X:)�6�bi�ڻ:�0z�X��:9�á�N���V���lB/�0
ee�>�}*�$��I�d
��U���Յ��^fC(���kK���w��`K��j~���*H�:}66n��6"+�Q�w�h�ifuIn�(�G�/�7 �a�ɡ�Z�B�}�2C�}��!3?=Gs�NG$�æ��L�#��&z�����db�8�g?��]b%h %ƈ�:���/�-�����85�n���`^�xW�9?$	��Htv -c I>ځ'�oy�y��-�٥�+�;���o�Œ Mt>�ÈQ��{b6����%�&r����R%J�#��$��
W(I�B�.��4(j��-�.�Y�T�i���d$���|E�A��1��: 89����F�Jޝ��*]W�{H�$�
������P�~2�G#��%.n���ѱ[|�X��HV�⤸\>�@U� {����]R�{ 9����%;&|���Y} �:��J�b��;��p����a��xl9����#e�8q2:ڻмg7���\��>�x;��<.������o��w�y^�����|���_]����E,�@�v�������m{�� ����#?k",�����m�*�D�ͮ�Z@������B�����>K�63 	�.�i�̒��p��Ɍ�W��qSq�#�b__�������EkW�<���[��s�GG����;�	C"��W�#�P4�1�����i�E}�ք)t��Ѫ$�ho�!�������(E
��mx�U�Jt]��2����d�Y�t=��G��G�>fh�����>�a�_!����%ig{�[U�k=�;B�V�2�Υ?EЕ��`atU����&q�/�F~�\G��	@E��@9�2=X��oQ��{?)7��<J(�2���0�U���<��>z���9]��xW��,ʃu&Տg�}�u��+������z^݃aÆ���M-{9��X�L6ǻ��JlU"�FΠBA�}��d��v�=�'�S�i�d��#N;�ˠy̫���u�w�uo�%I�弦cw؝�	f��j.�۹�	)3�\6��QcQ;l�_�.\� ��a������(vzHn�HѰ�y}�%�p�0e�tȭy��+���J�F���c��k��YՄ�2�m��M��	����<\�\�X�	����.��d��'�zQj=O����KCq:CѴ���=�(�Ѳ.2z����l�Ϡ�.� ��(#�fiZv�D���ʩgI�#�>d)���CVT�ޥ�:z�d"�lC�$c��@�&�5T�ق#�M�w nj$�婔�EAd6���L�8r��?d�OS��s[�������dҶ�h�y/Hzf��Ks�(�R��k���=��F&	U��kn�e<���0�+����>'M̭z������E>&˂��sq'���DfA�i�(#��!G:Y�"�	K�(P���͗}&qQ!���~#��X��)-��s
��t��9��c���`I&1�g�t�M@���O���b	��W��
��߾�t0��g��+��_ ��{@��ߟ��v`��]HY:
��dJu`��!X8�5Z�?^	?��K6�n���S��ȺCz��wny2�K9����Ƶ"�΂W}�)xe���__�D�ˆzC�#!��;a����eh�$��>���s���������I��67��mw݃���=:�L�%.�^�I��`��,��o��9������{q��7�����d���/�o�u*t�bj]���G���W��ԀX�9���؀�\�C$���c�ct���d�?m�A�?�t��GC\��ܸ�����L*sL�O�m�_z��9��R36��C�/*S.�kű��{��
� 8���;�xҀ$k(Xy���-� �@<��C5�,��ю��S8��'�V�ğ��&`S^{�%��t8fro���i��b`�-�6�P�,i�C=��ig^Q�ٙ_��$�`���m�ɸ\�>�M��&9���Y�f�hW]C�$:\P��I�`"5�A���"m0I�O��-���̘�.|�� %�`�Έ��O�4,:�b7���F����v�_��J�2ȯ�@%���r7������R����փv�IU`C��e:ޒ2d�NŇ_Skiq��ԐM�9�6l����L�T4�,?��*���N2E��]vn�࡝�9����)�+*�pѸ�4��FB@b�]-���چ
#��hbzmba
<���"��ш����BxA�D��9��?�� ��ˆ,����p�e��Ԑ�t��&�]'�(4�����z�v	��{mJ���<����#������@�J#���P�����,�A#GGEE9�^�KX��jC�"�Y$Rv�nB<����	Y0L�HT(��Lt�&��%���~)#�dڀ���8��bS���$eqޕ��J���QX�y��b})񋀔l��]�~��8|�8�%��a3>J����<�����!�>;�0x��+���]�"��r/1 Y�� ��5����� 	�e�V掮�Q��1�߉���BXQ!Y9R2��+ŉ_�/x��>d�Y_O�(��l�t�@S�flۼ��ir<`��yه��w��Fљu����ҕEo?�k�X�{
�_��J�O3��e^�}�/Q�8�b���~7��;�G�%����ظ.	�d!��7�q�O���0[jNfE6o�M�����2($����',���*ܒ��ƆV\��.t%i'��E�XP,i"V�a��@� ���\�T,:[O%L��!��u�E����E����K�B�� ��x�g b;�94��,~��^��	���{�%�Y^��ϩ�U�{rI��HB$0Ka�%�����m�]�����l9^c�%���Pif4A�cO��|����W���Fиk�Y3�]�������0�sW�jON�ٙ�?�ѵh�h����
))Q�F�|[����B�<������MC�Q�N#}��~r//��k��G�~N0h}��m/�MD����̢�A��D�B��x����xҕ�xFN���"�*tjuh^��4��#�NQ�����Ȩ�Uĺ��n8=�Nd"bX^	�e��h�t]�sp�!��b�J:'L��n�(Q̷f�)&��8뼳q���Z��/��#�+���Aڽ2->Q���i<��VB��z���Y(�T'l6��r����Ix�����8��O�t_�Mlc���8�SY�T%����k	H��"��:I��p�P�s��ѡA1-�9.�97P�c��q�ˉu1�iXr.�+d�N� *�C*��"������[u�Ւ�3-r�����-%���H�����( C����G�h#�ZȂ&�����rl9k[�ߪ�1���V�\*�6-������F=H��c ��L=�}�-�rr2������tuN(�߹�>X�L�$�<�Σ��H5i�G�������ܯ3�6�tɲ���� ���:3H:�M�ҳ�y�@r�H�O���������K�B!�,���ai��
<c���ܮ��/���dv�ړ�Q,��j����>�m'��5���b�d�x��Q\s�0V�px��0��`e��t�q��oD~�3�?{��L�[�� y�z�]�?*�A�T2� ��v���L�ٿS-�Q���D�6��2@��c�w`T���%-²�����ߗB^g��Y���}�����.�����E���a���h��ڗ��z�v`��Y����_��p����ld~�������6\�1�'x�����R
WY4���,f�pOb���ٿÚvt��eI���cں��9kd9�쟱~w��Q�xI*A��~b"����]� D����>�4DN�ய�$E�^��C�ڞi?;��k���!�t$�۶t�;.��%;�rq��9J�U���U�W,Cnd�����E�G�2��5�C�Ԥ�xʡ��~���!�2ĝ��P�+^r���S`�5�ښ� m,���/��6�?�&�38�����`(�O�´MU�r��=A2'62��B@��Ih�g9�(�NY�*���Ȑ��հ������!����)�&���X�z��&��$�&Hc�cX�<�ň��d$�K�W�d��VMD�I�:��$�!����D>�b��5x���E'��`R�� �y	��I�F���	����.��ɔ�.O��7Ě�`����-��KM�z��𐈼��	';\�V��T[X�i�L�Wo�%�g0��Q,���Y7�17='���o˱�D�]|�ӕJ�nT�	��ufe�����\����3��m8V
[���8F���e��q%V�0�_�ڵ�eBҨ�!��2]�q��R;B8��pBh��whqn�T�y9m+W�M �4F;017���}���@؉������ALZVf���,��!Z��y^Lc	�
���"JХE����N,S�8ee���$�%���td��p��q�����_~�9K5���z�CO�X�xN����?�xh�L\y89��v�v2|����'O`�M��̀��xΆ~��1��3��� *v������+ᅿ�+(o|�3v��۞i��"��������B�ڂJN5t��P�����7Նӿ
��%z�#u��C�wBx�%ڎ�E�� "�v��6�b������C��]�J����o?��w�\3F�	D�k3�+K�`�f�� 7���[^�w��ڞ�j�
X�9�~�-�3�BB��8Ī���~ꯑ�; H�����0j���t{e��0ffГ�4·>s�7�i;��g�^!k���7d�Q�|���7��_��m�������ww������`*���,q�a��"M���(]���Ƨ?�5%I��ͣJc�[w]fzt�Q���b3�ˮ���+	�R���H�>��~8���ŝ���+V�69�Fua�C
8>TTâ��?�gA���>�&j
�(D|/nG�t��[����6�_��}����?� ��QԘ���N�TS��8��!�b�)HBo1G*�AM
B�;aȥl;+?Z���֤�,#>&pS ̢�� �˘KC��)J�v�9Z12f?0�{q},C��T�t\r,�(�Rk٘��e����4�������}^M��ps2�������
Ĩ� 'Jt�Ru0u��@�YK�TQ���lG@R�y"��*}��uТ{٪�I��7�xHc��y��J���*<En����Q��FGe��t� �����#.R|)I�e��qۘ#����iș�qPք��/�eX=R�՗_�^t%�����]���4j�����sĎ�Ե^&��-����tw�xF�$���t�+E؟+Q��-[ ����	<��v�صS��\/�"�8q4F:j��F��M̴��L��ʰ]��
�i����I�u��K%�hJ�i��r3���x�ˮ���'l�� �]�D���}�.���x�
��r+��ç�
<�cW֍c�z��zRcVFߺ�	���!T�1�ƚt�/YWgbK����Q@�AJ��m\��Wb`�fhކg�Z�?�x��K��Yر�~8Hqh�t�]�燍��5�>6�Z䡭ъ�X�u��l�YXR�����x�C�[���b�L�Wo6�D�u��x�����q��D@{L�1�TC�pmZp�Cy���:���h�LR��\��7B+�´=D�.X5���ۀV
����/~��?B+����L tM�_-�vK�i��"|�+����`U3�7�j��ܖi� �I�eCE�����P�J���C��}��[��8h����ٽ7z"V�q`j)��,����ËV�ھ��l��S f�h%���"Ot�𓎣�*��D��rG��p}#�������h�L#Y�]:�h�nU�͔z[���f���,�H������]��'i%:��]�p�������������?�}�c@d���8)���Es0�x�{3��z���$,(E�, �6ƜD��Hl��^&)n�Jۊ�feLX<�q࿕� %��(G����4Q3�������+�~��K\�RI\�C���pK�5����<iS�?�x���1K-R�j�M�A�=]F��$�Rp�w���M[&R�(H7�.I*�O�m�lšAY�N��$f��U�b`��Bq��+4)�ϧu5�jB�Zv�������P,W�l�%���
��P7���8����̻P:S-�U<�>�݄i&Ȣ@2U<3�p)t�����S�3���o���2�3ۦ��Ȟ�ؿ��/-����\���jg�e�{�� ����5V(�b�j�u'� �Uq˒�s6 �C#�X�q�Ɩ��5��翌�v�����X�j3w�]�<f�!��]�B&gщuĺ�ג�K�%��$\�����/Mh�)���ˢ!'C\#��"�I���x��g�D�ᒋ6?#�����ti'�V�?X���g�YZ�Z��O�Ϛ�� �#��[�w�a �đ�(̐7�M\����o�r'��H~n&����u�s�z��(�����^o�G�eY҄kgȻ�g�Q�,?|@�]�c`a���b�����h&4��gژ�k#�l�O,.7,��F~d-R8l9D�C���g�9X��3�ګ�����v��IH�aX��-�i����3C���ͷ�a�&4��]��{�X�����^p���{~YӇ�z����_�νX��\�5;h6���gǜ�KGcn
����|��(�	�)���.��u�<�u|��?��찋��}ھZ��8|����Ħ�O����2#bnj�9�}��lh���'��7���;�]�����B��|���cM�ˬ�1"��*ڋ+�!-��G�#���Y�t���O�Q�OQ�RHb4�N�ޗ�A���x�2Dp�0��Sz)Xth��Mo�U���o�;����w�_�&4�,Ei 7nl�@S�p*�ZѼ(b�6z��%Ff�U�0`Iv50tTs��̍(��K�H����I�C����m��Vؐ����Yrs6[�킲��/ȹD����.d4�V�[`���~�����|�S@��9]���i�ݮ�>�ݪ��cc�q�9��o4���1{�0�b�X�a�f>	���JJ�L�Iv��� ��2I��`1�F&E�X����	����h貦p�`�PpF��?���Q�mN�؉c�8q9e�O���jJ����+G��d"�A���|NhCKM�L䄡G��O�]��6�x�����7��_�t�ص��~F��:�{i�}���qb�+��1x.�'�V4�p���O7�&�в���N�)ڐ��qI�����BŨ�k��m1�r�ƍ���cxl��W��w���ë����0و��rdb�X��� h@���׀�1�W�1O{Ӡ�]��#��uq��/ b����	��t���T@,����?т��݈��-����
<�g_�	C��� ��6��~�>��Ȓ	H׏EwQ2j�xm/=5ZG�b��`�I��"ډ����K���-�@�rS����Y6�r4D:q�0�����>���IT�2�!/z���8p���Fbb��c|�#)��@˘����%D&�!��aZ:찃|�����=*�B5�Y���Y�������\#bW�
�qHu4<�_��x	~붗#%f}�����嵝ڌL@>���D��VI��܁O�N���\K�W�8aA���Z    IDATOϰa�
\w���o�N�3S�H#[[�i{�,���ߔ�u)��n��*��k��v���
��Trځ0�������IL�΋ނV�,�n���x��.Ň�۫�]���WU�����g�����ъ�����q!�)��*����!.�P����89tisJ�M�C�:��)�7�p�|ROQ��s� G
��!��d����5Q���[`����y I�B_9�����������������w�m UJe#���V%��� A)`�t)�_)f�h�5�a����-gBw\4�m���G�H���L��~�du���nK�ؐJX���T1"�HR��2�����n4E NA���-������� �����N=d��qm4�J�^�
�֬���8{�Ah!C(!�{	�>�2)q�8���U�B��6t�M�s$�%Q𙢭���^�F&45���)�|^� *P���ĸ S��D��|���fci�CO3!���*DP�p��Vby�"�Q�'�(�D��I�c��Q��Obհ�;��߱��C�^���q�NN
X����Q�I�}��/��������2�kן;Wk�\����2���lvf
u^~q�A}a�3*C�m潘:֮_�gn��U�F����3��4N~��5�k�_�q|���U��>�� �n�֜i�q �Dl�{�;9�ic�L"��d���_�瞷Zky=���_�TC��|y/mǳn�.�g�![��gr~l{��$C��13r�u��v���n�6��	��u�iml�q�s�#�ڍb0�e��6tu�K���-�As`�~rncfwF����Hc�	�?���v�܉0�Q,Uk6v�?�#�T��z���صo�O.�x� DX&1�6C;5��0�}R|�qcE���b�b!&�ò�G�1|����2�[IbG5�D�h)���ʋ�o|5<��V]��/�ve��?�N#v�/}�oq��S����d���q�f�r�ݖ���en<׮��E05��t�f<�� ��������0�6�r>���P�AB�,H4�$á��w���GG�$Я:?��˗�s�`8ga��!\q���������#_�[��.sX�1����E3�S�� a�ZC�ʕHr9��@rK%��Ut@ڴ�%��'$�q�:�{z�E��^~��Ű�zE1l7��W��0�L��A��kWc����1���6HO�ͮ��=�E.��BЍ��F������EL��*ĉHe�j1)�qۡL9� ܸ� ����%ٚ���A�rd*@A8�ܩC�d	8}����$J�9 ``����.>��Ϡ22�F���G���uqy#Q�,е,Å睋��b�c�c��1�v�%}N�#�<q�E&�wC4��6�@�:1��_P+@��쮳@�:)g,SMn8��/-t	�R%xN�8Y���D�&\�^�zo���"��0��Ԑ���v���3���X2a^z�ǈ3�Hm����4Ns����l�8gc7\{^x�9�N��}�Ъ�aJ�ϰ� �Jh��/c������B�8 ��O��'�f�3�8��9�8h�լ���Mt .qtM;��s���-[�;��=<��::����J�W;�mg��5l�s�]A�r?!��؝ �$���H�&�pM�GU, $o&x�M���s7��̡�3�܋�����3�����K+��K���Yڮ��
�ࡇ3:`�~�
)v��X�)�`M6Y<E+`�)����7]�k���Xїa��H�,��\�g]��u�A��ޗsk�ɬ�\�%R�]3�m0币��	�~b�9�Z������6TC�7�NVBed|l/f�:R|��ς�V�¨!O�БBh�
������%�vŒ3����|��G�N,��gQHkJnA�Z��ė^s)��;�A}��b!�`�+_�<�����;������i��j#[7P��W�Lwl�+�� ���/��c�L-;g�,?���~-��7���6���j�,{��؋w����/��2��4m�ᩌE�y+��q�1;O��+��tx���t�U� ��`v�>�BeD��(f_lYU���oE_�CI5�n��j�Bu��0D���ܜ�4�!x�NS�����{�=Yab-N T���XdJ��B���*/8	�a��ᓠ-��-H�t���A�1�P,|��Dh���K��+����|�h����ʶQZ��i�1��$��ئ�+1K�h��jǆi�H�NR�}��'��o����.�b-�V	e-��o~#>��/��l�U�B9� lu�pR@�7:r�6�u124��J�ӳ8�c� t#	H$�������S�<L��� �4h��G�x�ҿ�F"b������$�+=	���(�`)��)�2�w��)m�LMxB��]M!w%=>�v0�R�K��Ҁ��䓒!�(��1P�ĥ��B�����U��m���1�o�s��>��堔�q�@;�Q������m>��/}F�hf67uǎ���I��::���؈�+�0�_��atjM��ࣸ�{�ɴ#�Jh�9�����Dm���"z�ap�KP�&��������!�^������e箅�Ϣ��p�yK����҇�+���8N�Zډ�R+���mY7Nd|Ҧ�L������#O?@�.���!�lŸp��k��?��l#��P�`8FW��[.A~p%4{͏u�5��ga��(l��R�z��B���m��i5q��!I�nuBĺ�zb��� ��~d� ��(|t7�<Î�b�l��m�Hm}##2�q\as#y���E�?�Bs����/��Gw��M%Ԍ)�	I��]�q4�a�_u9��G�E�&�C���{ٛ��+R\�Qg�,�K~7��uxZ&֮���桼�.�,
��p#Ϟ�JM���0@��0���d��?��������8�ݘ!v6��l\�_y�X�|�jڞ�FF��A��']q�H�H����+#�&ظ���W˾�/w�O�⯑���D�s��H%�R�(l���vW���K����B}�t��@U��D���P� 9VXG���m��$ t���>?�#�'9 q��$q�������3��1r�
�a*�zQe$�NWv�%�[�$$-�)q<�g�	�����tX&J˗�U.���x%��Le(,�ā�L�Q:&Q`&+��+����ĝ��XF~L�����+e�x�-��w�D�����)��{����AР5m,@G�����7�+��ˀmnE��%�P�d*�5攆�?/X�3�3��Z��Wt�2-Z�2|���aQA�Aj��P��@Dt%&"Rm{I�B�bN��I�JU����s"�v�%R
�� &�Vb�Lpõ7`ٜ����u��R	���(������u <@ÿ�y��M/�M/~\��c�`�c�\� ��0�Dk^��e�0�j�o��Ǻ�=�/��G���q�]��7�
��j0W=�y8��8l��>���`plo�MMr���c����Q����E���NCQ�,[�g����}ŋq�����{�O}���-�vi~�V`���y:K��3_�]����j��A�˴c�i<���uD\�J�vWR��0����'񆛮Ɛ� �qZkN��`�S v�rY�	W��e�tYJ������0{�ޤ���=a[:r���1u� �މ��e��h4;Ь��csm�1	�~T;�Z���}�&`�t�)l�d-+�l��QD:ӻ}�tPj��o��/{1ffObj���}�8<� ��#�n����qr�E�IM@��������pË�D���/����.4�N����x1���G7C]�lC�5���*�Ƚ��\+���yXWr�O��h���}[w��V�VFь�J�,8I�0��fϹh~�5��y�����SӔC�0[�g����8��>��O��8�8Ĳ�05� |z�f��Ĳ��������_���ŕͯL4��l)s!�.��!�f)��$͛���{|}ܨ���&�l��@�'O
K]��PeQK�����D�� �;0=&i'�;>r�>E���%Y[�=�C�腚��%�Wɏ	������PȮ��6����0�9�&(�Z.�&�%Z��vS����pW���*�X68�'�H2$�$�:(�4O0$���i�� ��2�3H$i��նh{���56�$g�P.�b�K����)5��) ��mq#��3��F��K���9G#1�y*E[@T϶Xܩz�Xp"B'��H��=O@��;v/tP��� ��qp�f�`�L�,���I�onk��<2�����9L�)�	t�CC矹���
g�����Cخ� �o4�Q��Ͻg�w!�џ����ǲɓ������k��l�[��Nc��5x����ə9|���05 v?R{�^�x��C�X���bjnhIL���Ll�-��핿��/��;��/���7��<�W`	�<���Ҷ��W�б����	4;>"̈́��a��ql�7����Q�(��M�L_�qfg7^{�,���	ԏ=��B��}
��:=�a��[_���!��#k$f��	E	cS��,Th7���j�-85 ���:��t�}	��y�������M��L7B<��8b�"NS�������GaZ9�<���B^%m��J1YA搷�#�h�L���(<��(Vqr����2tH3	"�nN& �\)����t���x�K^����kp�x�׿�בY}�S��a@�,��ޗ0R����9����v$Ȳ����dR߭�kB�"�5��?�9|���-����	aJ)�u)4	�+2��o�9?���ٌW��blٴ�����Q���	
9ئu'�M�����{T��S*�I�&8R�=���(����1Q\�����)>��c]��/���Q�r�.:����H�d/G�ŭX�
���j�"�Dĳ�t�!��6RqϢ=�
�[��6ѝI��	(�N3�^N�|�B?�j-9��IP�+� BPң�$���w.���"K�#��q�c�H91D('s*֪BEb�-l!&�����Z.'��mw`ۮ|&5CE��́ð<(v�	�[� ��*׮\�f��F�#V�+���,4�0`�����7�ol��y�ffН�|e	l�N�"�	>ݒ�;����!�~�X��QJM��Y����F=Ӏ�"
�NQ	>ȢW.Y`�9�y��G36:dC�"�7�;A�nC�9	D��&cVS�A:ߒs�X�Xr��咉J8g�0�XQ�U�m�u/�_��� �[�²�0S�`d�l>�\���ܟ�Z!��d{v<��Y��k$��:�(��|�r��Wn��������br.@7�S^�N�bבi��a�A7�Ď�r
2��a��4]�7�I���%x�s� B[��^r����Ŀ��pi��X�x��E]z�g�
91���B� &Bs0���][��#S�n����E%��I�*�l�Q��6.=s�F�0��X8���>�V��W~zexc+Wb��͒�̂fv�&���b	��I�*"S�!`�I�0i���p���9ؿ3ǥ�mX����*�{d���F��V�y���Gь��#�-t��]�	�A%�@\�H�a�o�".?l�P0�;OQ&]�RN�,tB��J�� ςG��J���ҽi,D0�z�
ٿ� L�0��lD���=��o~)�ܰJ�B�^�|�*4!>��V�� �a J5�;���b��XhFr�h"��R��5�i(X�	�D�	�`������C��kn�V���Q�*!۳�Pn��znU�� DJ�
����uzZID�;��E���h>*����(�h���W%��m��dy5u�z�ۤx]�ᖪ��-�~Fq�K��i�J]�/�=�W9�C�Ձ���Ҹ"7�`�6�\WZ�r�\�����w�;�nN~O����t��Ӿ�6�����np������z�3v���.W�;A�pTAM�����i�vt\
B�fDQ0Nѷ����D�n���T&I�K7ތ���=L=��+b}��>�{�ݘ��b~fQ��r<���+\�Ҙ���$��@xM��*�$�5J����;b?@z�J2�} A�W����X��	:�����Y���	�˄L@'ej���Ri�Y�,nöu�9]�	$l^;���a������\�����������v��y]�MϿ�YQ#L�~��]�A�Z�� ��,Z�:n}�r�,���S_�'DFs��VD`p�இw"ы���hS���u]y&1�i�<��7����Z(X%'�����X�g�7�Җ��+�t��Gwi���+p��l|j]ܚ� 51ۉ�/�Į�s��^���l~�%t�����E8o�
l�È#�?��l�E�dn�U���X�l%�8g�BF./�o��]& �6����`��05�u;h7��똚����<:~C�8��P7�v��ڊ�����2f�)��fh��x�ZV����\q�2
X�`c�B�������ҶS����c"�[B�"e�0=q�](;�1S
˰�k+E��S3���	\Oٕv�.���<�h�]��o ���ۜ<�"87�|�(�m,|��G�P���o34,膈S��y��%�,"U�\!"v��KĲWevH^\ [��Ժ�Ó�y��,�a�srh̷%���p����*ԌT6�Q7����,b� �R�)��g	R�bdt��2":�66m؈�B�sU��E��󒤞�8U�I]@�c�+m�,;/��Ч��T��$"S����ϖ����u�I���,C�TDDG/�Q���Q�Q䱠`����&]K��e�v��R�SX����P?"j�5~��@�gb����Ԩ��g����.SKkbFM>z�}��!�AS�U�4��bN!' ������E����?`��TV��K_�R<��CX�V�0;��`M(c<O�+s+����A� q*C�9��)�ۊ򾗿�<=���q�{.�I�)�p��� �ni<Ɗ�E� ?>��s����(�&pTM�R^?�'e����A�G��)�K�P�[H�Sx����Wo�}n� ��0Sf��(��aht#.��UϪ�`��_��=��&���y�10ߘ�eϿ�\r9ꡆw���04��U�t=B��������0�4:����=�2�a�l���z<��Mp��l���h��_BK/XZ��"+���9&K��3\����gSs��L& af��\�n?�mNb!���:t��md�t
jKҿG�r8k��0l���wc��Q�4s��tҩ��ox��$!]tQrܜ�7�h���$�f]\��;!��f��s�i�[���p���L#F��Њm�(��h:��P�A��u�HU��e ���]���T@@�+�/�Rđ$���fH�E��Sy��4z�� Q�̠���f:q^фXl�y&e7;C�U� v��8�<AAu^>� ��g&b��\//�¤�����Rl����"MQ�`�;����As��T��H�Ŝk�!,Dv��/��&�����Ύt���I"��B��*Ŭ��qf�IG$~6-f���N�ǅ�^�n���ĸL'F��p��aq#㴁 ��k?P��*��9#�Ɩ����I�-2-b]	�Sq��$�m�\�,GRD�K���!!��'}��dh�/����t��� ��r�Yصg���v�.��}h��2� d9��3�BszA��&��~Ě�ֈ�D@�����C�V��_�Q���Bf:L�g��a��"r���Q�ӺH^	�]�RY���]�s�9ľ=O��:3��3���eo+ڝT�4�y-鹢RIR��d	id���n`=r�v
���ż"�V
�кZ�`�SD��I�
�0
��e\3�Ҙ��',���kQ���샳�Akj�W�I�y�:���G��_ǣ~ǏDSw�RY����p�(������n��fvp�64fO �س�	,[�׼�l��9�����XE7u�凱���M�pr��n����:2C���\����B���ҳP@�E֬\��~Zw�sN�X�xN�C��COgv�ޛ��j���    IDAT���6����'g�Ю�غ�8��.�o���z�U�o���1�f�����V�Ɲ�r/D�mQˇ�S��D�טi���8b�+d�`�2uU���,R�����r ��nU��$�6��n��T�P��D'u�G.���g%�����6�p�T��l��2?�E��"��'_@�%�#i@�d��-%�lC�0JLOt۳��I��=��U�bZ���~(~��P��k���I�E]x9���Șu����b0c҆$��E�*�)eg�I����K$�(�(���' \Z�ܗ���3�����8FѵE+�v]&9�H��+L�gdJ�@ �|���½/�Ѷ�b`�R�kczz�����l$ٙ%C�k�D����9�q�3k��lE��er����|�0H圱�"�>�ͷc�̎|��J:B��Zb|�r��vS��|���pީ7`�׍.\�.���\^��>�8���AF"���p�0`2[&e �@d�!zN�lW�H0�gxR�-ֽ�>e�='R2�! ��1��ʐFN]�HK���Tz��խ'��y���m��y��J��4��}�֐s$��Bc"-��3�1M\�ȩ	�i��W ��A"?�M,TB�S��*LP]2㵲H���,q.��zF�c�t�	��VH�>�Qb�����M.	�z�Ft@�������5��QtSl\�;���uۍ��|�(0����a�E7>�k�xfW�0u��4�� U9yB��ӿ���w����̲�6B�N�c��q4#�ʘ��r*�ۥ���s�����3VÍ�X3:�5�G����t�/�^��Og�.���zK�=�V`��=Y��\�F��h�����<��j���B��x)��d�?
a��v�Ӂ�מYFu,��F+��	�JaR��K>fǞ�n��W��'2�`�����jpsy8���#�3��509�ı�:Z��@����щ4�:���eD�r����t��q$�F���|_�bY�����.��]e%�`A&,��g��N|/���R_F(z`a�+1=;��~Չ�! "bfK�E(������Ȗ@?ۖ�O)���^�ѳ9��E�ChC^���=8��#�����q'��E�)�{V��d%<$����jql]�p����'5k@�#f&�]��P���+�b��w��5��I��b��.�;���qt��r�=87�m��s0��W�''&11=�����j�r4�M��+�)]���$�,��:�	�Ȅ��1�y���6?���F�s�99�����B�9O�9^em���$A����E���ӁJ�%���%��z�$ֱl����!�H�N�$��/:76���?)��e{b���Ϣ�;Ć=��mJ��t��M�FD���*;����c�a'@�)�r�(p̃�/�����w
уI�W����C\�d��m�H�7�Kae��1Ӏ=0�& ���3[]�C���~9S�7y� ��_ߣ`Q#S�}�w���)��d]���3�7��z��Io%o�YN�=C}��8��_r1~��K�;ޅ5��+�����UV��nDa�ٟk�̂���;��v��|1�Gۊ7��-X��|��{q���M
���%,D6x�(�υb�A��iy�ekr^�ʗ��c0�l\1�@N�
`i�~�+�@~����Y?�+���=Y�9��n�a��c���C{�IH=���#����1,���G�Jf�B�D$Z6\��ˋ:*�+n�`���tQtD��$��5>ؙ^��H���������4�TTx�f"W,c��đ�,t34#� �J��6�	j���uh�Ig�p��QK�őH%9�͗g:�~W�Nb*E�v�����J���K�4qzR�
�%�AhA*P��G��1ǀ�jb�.A��^�G+L�+h�����C�̍�9АbͰt	$3u[
�DOэ#�Mh�#c���:�T�8�d���r�Z����e(�'��pt72����U^=6����Й�P�cC3)X�ʝİ��}����@_�t��A������q������O�<��\�F��Į��;P*����	<�{9�rQ�`ddL ��ǟ���:�v� /?��j̢�&GR��+��z���9��W�d��WD�:���A�a���))z7o�,%q��Q�</���!T*����D���{LM�IR\|%��$�]j�<��p�y���M9�b~G��$oElm	Dc�4):���R��sU�Fl���h@H��%�P�Ç���LB���@C���-z7�-Q��x�,�D	C���<�q'����)0��&�kq"G�7���S��� �bN�Lz���]��I�����
��QW�2^+�l�g�Z�ɜi������Ll��8B��!oX=l��]�߸�ztf��_��e�^�W��/ǲ�_p������]���};0{�*G�������"W��7��M� b��4�Cs�4�j]��GlXȹ&�,@��⍷�.޼F Ț�A�_1|ڬ�������v+�t�v�ti���
l߽7k�;
�8A���t���vD=��ư/��H`��E.H7a7KZ3�`mEǦ�
J,�� N63��3�)�0@G	�`�;�a�U|�,{V��6���h��g�O�d��*��PC���\��Ԛ1���Ff#Mu��D1�m�퀱Ҡ����k�z�ZmT�<lW�����ͼ,/;���RYRL������)ɫP#:+	=��⸔������A�^��%�+�ت�͊2�
73�"@6R��%ޱl:�1`/F��⤤:�tv�ى�.n��6�To	^ԩ��aOT�^��E��p���(:3�H)X���nL̃���QK1:X��^v!6�_���<�֨)f�g0]|��x��W�����o�s�!��d�4���e(���nX;���}���Z�#2,����T�n�\�"-�����]�믽��6�}yl�k������xx٘�ף>�~�q�[ؿ���/�A\�d=i���=LP*�P.��v�_����~[��{�C�ބmq�5��{؁����ׇ-mMZ�Aqliw1�)l7/.C��c1�OvɦV)��s�yp5��rJP�C�.8��?���!��yQ���o\qc�|ҷ2 O@N;bS��s����)b���
H�& 2!1��*G,��)�" �M1�� ��"���|�����s��;j
*�*BNKdr%���+A/�h)�9���y�f0Z�r��%Xh�i��H���>�W����m�C�n�k�|?�y�a&��s.y*g_sZ�����o�"��qd�8����Y���>�Mg������:Qſ|�̵Sh�L�4t�A|硽�m����d;�w�Y˃�7����հ:u���3O�5{:ߛK�]Z�g�.�gՖ^sڮ��O��ڊ&@3���`��=��ɨ>��
E:E�J$+ԝE{M�X�H��1ʮ��r#�6F�8h#��C��}y������|��J�.��.6�d��l	:~�V�Y��Flx�f&f[f�>���V�4d���"L��%-��-)�I����Q��D|쇑�RI�C��K�8�Ws��9��E�@�Siܪ�z�wJd���e�|H	Pȃ�!��m��B�"���N2��)�PB.v�{�N3�D� �)EU� �S<}>eQW�rP~�(��'���9눙�Єtae�f�C ���E��5��y~�u�����(?�������b�m9�G�ѿ�'��}�8|X��y]�������	`�unب�7�t;n{�/b���{����X�\{��dv��^��W�
�hw:��jx�/C_չi�{��K6o������ܑ��]wa�����W����H�*N�H
�0�J�{�%Nxb���H�b�K���E;��j�s�t\�n�Up��m�-9͔d���yO����/fʐ�(�8	�P�^�r�)M������i@�"�'N�GtVԩp�y.~[M�����f=헮#
|��p[n�(�s���ב��d�m�a�@��eZ�����-I���8����=����-�R��}��'���5%�՜��5%�,e����@��7��èU'02�L4;+7������Ӷ8���isS�X��䉣��?}o|ݯ�y7���f��}ni�ā^^��'�����,� �]4:>*}�i��q���[*8K"�ӶXڱ��
��7����-}��;w���A �m9�2a���܅{��GG�#d��N4B�Q:)z��A)�U�S[Q�4��c�b#ge(�ܤ��Q�N�K&�p�V%-[��qA��za@�\ɻ�x�k���P�G�"%a�����w��H��ud���4ρ[*�+����/���8>X�	��,�~���w�g�����c��GܳmF�w�H1�HYa�H�:'*�"H���%!���t@H_YoS�m��T�}yHz�nR�R�KG)�0I��m׿sG$�r�1Z3�@�����δa�tł�H0:�Ǉ����x���q��lͺ�����[�w�m۶���	��Ϲ�ؾ�I��~7�cڟ����ފ�~��p㏼���z613�1q��~�-��E	��.
k+����ǎNd�^|����C���#��.n{�o�����;y��2]�Jy�}���h��tpb�!������jyl�>�	��,��
Bδql�A���*̱T��n+ay�y%Z&�se�۳��e���!�w��n1wd1�]$$A6ӱy�k�9-��y��4�F$� Q��_�
0����
�Z��W)��33��K�:��hAO`2��1q�u8�g7jǦ�k԰X�:aW(������D0R�n�a�X���ؾU�����{_��L�l����8��+�-����NڞEq97#�pt�T''Q��Úu�q�ނ?���r+����y��z|��'ql&��VD�����}����V"�Y�P���M�>����[{i���+pZ�|��ei�v+�������PB'�����N���!�2�f+~N@X��J"���
%����1MG(%iL�J�����R��@���&�K<K����D�2�膃$#>C��fw���F�F;D����	S�,j�Z�#����KSqۡ>�i��#+����Bc������lu{�����T��by����C�D)M��Vӛ�p��L>S�z����o��0Q��dH�d|���� ���Ǟ�p�@����(�w� ȩ���G�G�j�/�"X�A�+;�q�I�R��`y�9gmZ�����q�������ĉ�ٲ��������;v�COfظ�0;����	L��P�+a�ex����e�o��7��G���}{�c�m���.P�`xp�{Aw�~��g��}�l���x 3|���(�p�-���>�m�-�4��|��̾2Bj��������!�E� �u��)j�u�V�˔�A�gm؄��<rASѓ:d���7Ak�����-��A��/�"���eZAZ�LAHݳ�j�ȕ08�^�$��uZ<�l���j��^��p-]8j��j �p�S��\Y/9R)L[���?{w���}a2U���&�f��)�;h��!�]�ցgrjc���e�������?��Q�W(�r��ף���������3�x�<3�7K�:,��4\��G�Ǒ���u#��^y�K1��������0B{���32s�#���{�u�h��V9[�,Ѱ~�#����X�S,���
,���x�Y;J�')"�8:[�w�>)B�v�G@�0���tOIߐ�:E'Q�N%%�D��$�:�md�l}y'�P�C��$��6�t�9�g̶  �i $��펏F����z��bf
h�>9�CR�{2YU�p{LXł��0�AWtB��J���<�#գ�,r���'�bK�~����%n��Rf��8�����?��C�n'��\Y{MY�J-��k��1a�_Q����sĲ���.���󅞕�p�	�D���Q�C+����S��nׇ�����k��W߄�>����;~d/%��MKQ,�)�f`��� �񓇳/����T(�V�� ͰQo821	ӲP�y�9���=��]��
�M�Ƨ��&fp���؍��E�,�n�h�0����,�W��{��l�:������(I��ܯru��i�l�AZ�$J�D2�`&��x�$?c�D��gc�36`@��q��ygf��Ω�}��o���"l���n����Pu�V����O��o��+�h��_p=�s�vē=p�����0�p�#@�+�4`���O��$I��9tl���%�YM�׬E²�V�8r� �b	�M�#!�0��������[���f%uZH�!�g+}<�?�� �6��[�K��z2�#���/α3͍���{C�7�IV�*�l2W�yw,�^E�'��hD��e����rah� |�Ec���q��!�/E�E�Ŗ�l#͙*_h#�57$t�(⶷݂U�6�?� ����ZIX�n�����3��g��a��.ѬN�P��<y�v<����F)4-��ۿ���=8zz��+1�00]K�=�1�wa%;�*���7��ضr fyS`��v��}~����n�7���!n�m�ؽO����ȕ��G��!	@�\�d��@�BbPA��_����Z���\�e��ET4���N�H�ɎW6%��ۤ�ʱ��I�	���!Z���5Q%�*Oz��
p*�x՗�.����
ZÆO���fjh8!d��Z��Ht.9f���_�� ��De�f�y�rkZ֖g.7� � 
Ys6	�PdAF9"��J�n	tI�L �|i�ʶ����,:[b_Y`��.W�Qǣ��I�jm[�v�cB�B��6w@�Aֶ�4�;|H�9#,=�U�m�������������ԩQ�I�R�B�s?��̊'Xd��\�)�
�+5$�q��%β����,rX4$i[ǦgH�������G�bq+�PFg�D�\�t� �Аsk��w��C��uX�Qu`��D<P1�7��g�L0 ��C�?���_��l�^�'��B�$�*gÐ�N $��Kְ�BFH;�ǐ�K&z�����~�I�u+�=�7�]��D���;rTf�P��"��<��bR�!�A"=P��#�FS��;�3�*ٙ��M�-��P,P)α΂�bƘ�ר5َ�锨��6��Ū((x[Ⱦ�����'
2R#���XS�~�*�܏��qΣ�T����"
%�g1�b��|!���QG��a�.��ގ��u$(���BK�`��c���������R͏���1�n�_��=;��M��:����������{����Y�D���qb��r�L-b0�o~�M�p�"��i ������?�v�_�����O���o��8���Bt��:!N嫸���xl�q�D�@cӰ\TG �s�� �ғYXkX2��U�3͝���FB#�JZy%J9�0o\�5�
x*�Z!nJT��x9��%{Z*����B' +�@�L1g�d
�t�P�WJ0�<v�"+i��$�6)ߡ�r�B.=k/Z�g��� �5���|N���*r$8g D���͈���N��(_��P�d�������Qxleu@�[Υ`�6( �Eo�I#Z���n©��0[���@g&��_p��:�?��ǎ@�lۼ������_�����w�0u���+���F��J��Ύ��R�K�1O8��I�^��P�u��_$�&`J5�T�?�T*0���iHR&I3�`-V�(7���ѴT8qe��.Qq�Oj��62���\^��M��b��3`j׮]��:���~��+W�����gψ� an���$��64J��V�O ���ZpG$��Q��4L�˧s��)e,��d2(�'V�\��l�?�8���t��Mn<�yzPg�� @ΩaO:{�D�QҢ��b��	�X�����3�U,��\���N;q?�4S )/�rr���ΩCJ:��u�t���$ �� ��C.p�G�1��Z��m!7��Λ    IDAT1NAe��y��ɂ��&�2
�Ԡ�&bj�i��,��/f�4��7_B6�D<ӃUۮĲ�?�u��'v����������Ӹ��B���z�p�-�]D�=53G�TI��=9�&����y.�8��CgL��M�5�xGm��=�<퓧=3�#�`F����*�T_a��O�ä	m�|U�`Q���j�A�d�Iu;d���\dH���ל����AV�d���i���&�����F+�����O���!S���F �(�ő��O�u<T.k��Y�:���ϝ;K�"Q'��ΝI�Z(�B�W��P�x��ӡ���V�$��9!�����{�&Ӯ�oV,΁���Cu)u"��(xP���|�ܾ�\���ʴ��4%���?*��A�i��SƋP2u�a���x�+nAw_?F®���(�/���]�>������xs�ih�����Tl���HIJW���aJ bƘ�C(�Gf�����w��1ʴ���ܰ8�B�i�D��Q��Oc��G��!��5t�;�Ju�Rx�N:��XK��~Ù��=����b���oa�g =�}��w��Cǧ1Q7 ��ܝZ��Y� �A�(t��g\��ٚ� ��r�&w�뺆��@5���&�s�3\�~�7ۉ�e#��!w�4W`d�.�Ŧs�5g[ �N2�~�s�A���=���Ů�c���x��`�����a�V�t.�#;�b������#�������&��<�LM��j��:GB"�I�m#'�{��7�8ɶL��MNr�b�.>l���9��%ӉLX>h`��c������q�w�չ)��x�Xs�۞���Ӈ�zP�
l����ƾ}�00�7��\��}��(6�J��F&j�q��u2����߸o^���`GkV��z��͵=���#��'E{�i�<"r�"B
��M=�骋>q �<��B�
����%�u+<���@@�zT�K�t#�xpG�����G@��' �ԔP�ղ�eY�Z�U-1��3�H�" 
�\����t*��v��BJѪI��>T�Ѩ7P���u�� �HS,�.-p��n?D-9���9�Y8����>���$��Sv� � �T��D�Xs���]r)����㤻iQ��!�����u��������$��`���N\�
3��Q."�W��N�
@�1n@�m���b��a�rX�r��ƛ���z���n�fe�S�� p8�b67�yv���fz8�'��O���AR�Gvf������'h���oxJ����ܴ/
�p(zuԴGN�b�ƍ6��7]ت��T��(��0�;��/����ؽ�(4�سgV/C"�B�1U��ٿ�&&�.�N��+
�T��pKD�#]C��&�'�V�m�L�"�u���d�jU�p���i�����>�NEf���CD�/$N$������xRWӎ#��D����}]��)��}�pŅk����,��(��&��_�*؉N�]r�#�!���B���З�L�QQ�'=,C��5��.�ܨ940���it|�t�ȦQ������r�4E�ꕑ5g�q8������Ӫ������]��[.F��=o��3'w
�:���C�:v���G�R�֭�c�ڵ�,�p�#;`f��7{0[5����i2�ݫn�E��A��biOV/}ގg��h��v�'�v��N���}���\B5���ci�L�ᾝ#x��Iu����  ���ЩȠ�|*O�6���%�ZQ��tRK%bD�� g-�89�ኩZ,P�ҞI���#��E�O�B�����/*�)lM��E"�g:����{�.#=��wG�j���Վ�ɥ��1��;���K�QA���nv<�<�N*h=t� ��)�� =Wz�ԂD?[ h^���~X��Xؕ��C���E5S�+���z� ]���) O��7���c�۴��t-��l\y�yX?��V�㧏��E����O�z�̀�Q���܇��x���I��	�CF4�frǃ��W�*�U�ܦ\rR2౴�&����	]TB%����^t�eН ^���ބ��^�GF�ctt�V������I�c�>Qm6�v�泅�[_����M��BԫU.�=�� �GK���RŬkZ�P7�6L,\��@�Tf�z�^c��b���8��g�(�@OW7R��������9�q7��Ϛ�D1�`Y:w����$��O���'���q���ݿ�\1��ѩ�����]I�`%�����ã�h*q�ԕ�S(��Pqv��)?��O�)C:)���=C����(#a+H�f�'a�qt��#����t����^���D�)|^��f�̉)UX�n{����݀���&��܎��E�z�UX��|h��_צ��A175Ci�֚0� �v��ȡ�X�d	�W���U+�O߽5��� �A�����$j��[_�R\�y%,���~2�9uCl�L{~�#� ���m��o��2 �5�v��������i<y��< !&��0_�
}.��ei%���)Wl��Ƕ,�h���MT�z0?f^̭E#r�o��!c�H+r�q� �G$e(�tQx!98Q�  n ���X����|N��Y.W�!z}k?�	�HtqV�D�-��e�B.�*�9I�!
�a��w�����"Sw�߀PW1>3��.�,Ugh^<��D&���~�� �cWZ�(����r@��@Nf��"�r�Jp�_*� ��tӵ���pٶ�HX ��J����c����	���54ƉHf���L�s}^@�C��p�l�|�	�H�d��l�1��%�6���C��$�Y�오r�ST����Ӹz�E��Z�Ge� :��p���;���7���^5j�nQk�qե���>-���&����R���iq2}��|h(� 3�h�.Τ{����#�щ��֠��c���������2�#a;� 0u���1�*Ǎ�I2��e#-ݥ$hgZ�P9�^�0���)�yj���Aa�4n��b����~y�fMetrZ����cӢP�!�ك�#'���}�����LŅ�S�s� ���"�.�R�?�J��T��L��+/���^�رG������.��iL����(gj�4"��Ƅ�b��1�MK������_�ʗ133��[.�e/�	�.{����[袊����rSx��G��ݍL6�ˮ1~�q�?��չ%��B����015�W��&\�a%l���lk��s@�}w�����������r ����1c'O��|ӹ9�	3с�#'��T��F)��B �5D�
Z�YxӪ,�B�eSf
p�E2S�Z�n�s�bs�G�V��z��U[*�%�Hrʩk�C��H��T�L���d�
iӄ�Jp! 8@ǿN�f��%�D���?*�P�t0�;T䪵�V� ���g�|����K"p6��0��q���d�oX���/�[o�Ё�<tֹ��%7a��R���0��c1:	���8��PD>"����&��ُV���O��8 �T���z�ZCج��qv_"���JF�B�Pp������7�W_��T�9 v���ZUS`�*�����n��q�kU�9������C�R{�r'�˯�=,M��z�ʔ�Z�A@�� Q(��PPT=�N!_.aq�a��3�Q��cvf��*.��l���Au������8���A�;���6�Z��	���W!4;��)�H��$�(�D&8�#��V����#�E��ȝ<�*0{z�NN#�|�\u%NM��ĉh�kL��l@��	uE����ey���˲"�؜���Q�74�dkM�{����8�,��e��K���)��6�d&Jk.�,3���O��|<�"�@���Ō���gp(��X�]��j��x9>��ތ�N�;`�������e=��C��8����0�	#mXwwf��1���1�/�]��ҕ��O�z	�����k���W���dC��>��
bF��xMÏ~x7���,��q��W�+_�.D�E߆ݵO���-7߈^~!�f�Cc/ذ�=�����V<G�}�<Z{�y#@ �Tk`|j5/D,݉}'�����>|
ea�5/ �y��z�59�^�g+%�EW��F�� �UD���x����K�������ŵq�%S�=Φ`�{d-ʶ���͕ ;�&Q3-���g�^�`*������bmaHˮ��A2㤥�xf r���(h+��?C�"�D+ڔ�-��֬^��h�V�����X�v=6nބ��ĎݻPw\x�É朘�!R�/W�i_�=Έ��֨< ��|�By�8�FN���R��ʌ*���id�&��ͫ�]o}=^t忟2qbL�s|\�z�	��Z���~$�Iv���	�xap�� ��\��0uH��8��s��먭B	䶍�TP4B�ʟD�w�-L�E�i�Z�|��a�Ƴ���1Q�p��qNI�%M�m�Z�������E��d�g�l0&$g+�&M�^�h4]����Ӄ���Q���ĉS���h4qᥗ`x�
<��v�OMrO ��#�}��ǊrTX�H0��|���h(�Sj�X���0�J��jS��x���/{�[ӃuE�rVlX����c��b�@�26[Z���R��{F|����w�} J��10
�����&�!�D��-���W_����p���
�U���Q%�S�w�~.�i<5���� �HXp�5dS6��)<�O�J#��7�3f!�;�[~��i����1v�q�{XF��,z�i<pｨ��fR�b�}�K��G���]�~�.�������n~	��d,���l]��]C��n��O~��@��y�����|#p��q���
E�3�S��y� v�Lq�h���<
McQ��V�Z���i�H��A4�(_�E gr�u}�%�nu@Z�?���n�B=:��dlP��&��RfBKġj�Lv;dI>��'F]���I葈;>�Ƿ� L������s �&�Jw��,?"wG?�u�$�$ʅt�bKc�����|x���q��!��
���*�<wv(�D��QG���
u�X�(X�m�yp��Ӹ��QWg�e�EZ @��u�T���tx,+�'�3���	Z������/ëo>[�}�l<9zD,Y�����O}D��j�@7�/Fw_���=5�0R�n����B�Υ�*��V+ӧ����)�:y�Wt׬�� �N�������Tm`��1�N�������o$�r7h8��k�3p�����b���H��(U+|�H�rj�4r�
EA������U�B���Ngx��{)���s��#Aȓ:��U��l/���Y�{v��]w݅U+W�\�����~$�0tC2ꨩ�]!��fZ\/�c�OE�~d����QfMԉ1���	v�-)K�W+�ozn}�EP`8�(ǧ�b�/�==�r���!4��]ʁS�BPX�E�1߿'>�'����A- 2�י��4i��Yx�<~i�y���޷�� �39f��G�ӳ䀖���)vʪ���2�1�R+��"lV��Nc�=����8yx�(�Cx�{�l��o��>Q)��К��tgq��w#?>���NT�%�����G�c����X�*Ҩ����7�7ހk���Ѕ��qᖟ=l���_�����/L��c��ßc�>"�~�!@|����ލ]�(�
"d�[@'����,���g7+��`*ӝ�H�nV�n���c�@�	�ɑ�a�'�{��V���E+�>T�"��-	'X��Ju���0m^��f��%*
���ak~l"��Ҥ,�^
Xkɫ�ܘl[���I ��	BX�"�O^��m��dI۠�v�/�O%y�ڡl�(����,2C��H��$+E�P��5 ��̔��
 a�����R������(p�!��(3��%�j�b�~��oê�]?�{��}_�KsX�z~��d�ٞ��Y����lAk�$J'�&ʀ��h@~3Q�TvA"����$w'h�)l�C<�A2��`CA!"� �t��Si�g*��L�5�B	CC�a$��nN��j��f��G�V�\9�L&�����1>�C�RE�T�jv`�J],�İ 
��e���<E ��I�Y�J����E��r�
N;'�U<��t>���,�u"�f:�Q�u�Z�8H����TH���D{�x�7H�N�Ǣ�$I�
��`��A�NC8%��b��Ÿ�GUFg��D�k�M�:����';oб�;��(
ҡT�x4��$����7�w7r�&�L\(p�D�B�Ay��;����͸�]���
�\0ܧ����7�{���<&'K����d�����Gɘ�ڑ����q�y��м:|M�ٿ���������Z��㇡�Cu���� �s?�f�L�ׯ�d���b+6�d�G]�ŷ� ���
\s���Y0� �W�h���qm��=G�}��C{��ރ�D�RC��Q�����O�î�)<SJ���a!9[�F��P��{Q���.�NI�7�,�4��X!�։�Z�g���������0��k�H'�ҎP��X��@�L�o�: x��R�LS?ӽ�_[���� �H`� ��`�K%?��Vr�# Ҳ�%*1c��J�h��&�.Z'�A"lU���R��*Z����� �,i���Q"mDk;�֪,Ԁ�xE���Ю�\��@`!����1' B�DUa�q�kX���\w9���Wb���k�ȑ��\��~��z�>L��@__/:�i��L@74��wax�2^��-S��[@ �lw[�:e�9A��98}�4L]ej�)��4��D�m��9#��F�Z+�b�&�bՙ9��@gO/�x��N��@腰�$���v!�D�����J��"#��G��C��l,��*aC�d��e�: l��Q8g2�F:�bk]6UP)��u�C*5��ј�q�����[�y�#%����P�<)�B97
�{��W�_?�>�����05�2	���iAs)�����B��5�����K�`EJQ�քajPM���b��}�x��}PcY�L�S4���d-��í��.Z����m�i�����X�Q���������G�N#����'�ѕ��W]�X����i�ڱ�]i,J8���_�}}	] 4,dWlċ_{{�>��?r�~�%�Z��W����afb]�).B����D��5�{1�E'�yp;֯ی�.��:2N۶���D{~�h_�~ёk��99�S�<\�O5px"�!�O�@ы: $f������ym��Ɇ7|{.�
��~%T,Q��u⇻PI\�A�r���[���y��D?��1�+�p>�,�ը���H�ZUa B.BT��%yv0��3�t��@��˟5+�08��E4��z�@���F�g'z�m:�Z�r,�r�%����0�e�T$�7w?��5�.�qam&_ew�l���L*�gf@��@%4�[Aa�*4���4n��
��-��p˨�J2p��	6&''y��3b��j����'�X��w#ә�a�������S� ��&�qN����B��a��[)K�W�0==�lH@ۗ�.���s��'�B���j��id(������6%������eÅ���f�({M�Ti1���3�DU,���1J�T���LR>�Ú��-:�4'H�""�u"���3��W*�wڎz���o0e�9w�����q�4F�6�"tݚ?�TC��$�A�� P*n�Y��ko�/��
�^�Eab鸉M����|Y��L+���ע���;��rY�����_�
��9��|�\��O���P,����D�*���+��;?���@���Fۢ����� �7^u	��o�Ө�q+��86�e���ow�O��K_�2��/Ǧ���m_^|��w����x�U[p�����#m#E!�k�a�ůh�����cۅӘ�p���3���1<��c���n|�+���;Q�	��H,�x�������CR�C���oS����@{�~%#о0�J�Ά�    IDAT��%ϖ8xhD���hP�i�
�Lp�Ӈ������@7숓/W��Z��8H].���"�[��L�׮����X*�{���\�h���t���-���6%��'�}�F M����Ag�Dm ν&�+�6�S�Ľ��_r���/���2/<�P���h(�x����]H��D-{[��Vf�����NRl�%;4�8���,�9�	Ѻq������G�E�+$��~�WD�xj�V����WG l��e��&�O�KTJ
�]-3�\�T�w1�x%m�9��u�P�#g���q80�1] ����׼���[x��< ��2&�
��D �s����d��]�v0�k`�X�-@���S��ا��tu�?����@E��0��K�'�ؐ-�n!fC��1|�̕��T(�E��I�}`����{!4��d=:��L��a�I�#˂�L|��Civ��u'���A�@�1�Lp�Ph��d�@�Bt�0���f�W�C'W(���:T˒4�փ�!�ܜ?�Q�_�K����ts�/�%+���T�q����m���7�NՑ� ���;ÿ�s�����~����7.Q��y�y.���+G*���g���~�n���>��.ނ�I	���H�˚xt���G>���d��l
�3�\���t"�"��3x�;~/�fkP��.�Qv��-��E	e�ɢ�+�����8�g4��7�r%��,����t/Z��/E襁����On|�(ύS�(44�I�P��œ�<���$b�n��f<�g?J�Wey~g3����`�_�0�eݦv�l������n�'ϯ�!io����wH�u��t���/p2W����HU$P��~͇K\b5�� ��1Br�"�*UA�:�~�@:a�&�!RI��B1:6LE i�8�Cf�L)W+��>Ҩ��6}���"5)�� %��3` z�L�f�uK�P6�1�	���J6�� <~/_"�,�pM'/��RYL��c�w�:+%�)"ש���ꄨ�|H���u�h�<�Z� i�yĖ��2O��─W�9iM*^���m�
�7�����J `��� YS�K��^(����R{%��Ô��sb��w����?x� ��Ra�;�J�)@�|���cp��|�B])t�t����XQ*���n���7J	H�q�������d�K�F�b�FBer�r��;�|�ۘE=h��~r�za(��Zi�VuLNN���('iz�J�ld�3�k:>�����Ê��
BO��H���܉2l��d b$;��A	�����d��-0�u9�Ç�E��c+_2O��m��%�Y�0Es:TT�h \�:RhV��Ul\1�7��e�ᚋ`���R�v&�r���l�>�(|�a|���5kz�cssbYW�2R��f���/�9����p�����E�m�괮�=>! fzz1[m������u��Z�ଡP��t�CdI�>��T����/\,O�}'&�ƥgݫG�B<��c���T���]���W w�Q$4V<M�h�x:����S�)��;	Cq�$l���?�0�O� �I�ҫ����(�:�d��#։�$�i��GҊa�9Nq�����w�G��6m �l;b��������{���[q<4���r�>y��?�⨻yd�JԜV �\����TP3-D��&������7Rt�s�H'����םf�I�&Z���Z5'���p]����� �J�O���2�$|�fe�?�R� %��:L��U�Ț5�z�:!\�G�҂HjV@�J�/_�s��dF�i�g~?��W
�i�h��5(ѿ�o��- e��w��9^���H º�����luIRR6Y�r���MNKl# Mȼ�F�ԫ�O4����N�!<�pK�ćo�mo�E!���cp�u�S�M�^s�y�cҖ���D��ln�L�h��}$RI�T����x.kd�����F$C�0W�c�t dkKv���33�N�  ՗E1���)x��7S��;��k ��F2���p`�~سq��`� �S���n�TW�n��z'��:��B;U=�rŀ�K�U'=�%��b�p�F�ƻ�wS��EZ��H�A4<:�t��2a��������w�(d0��Q��n(�e4cX�p�X?����iY?V�%��=��l�� �<�0��A�<=���n��?����$w�w�(>��#;�P��jQ���[��oQF�kbE_BvVf�buOZ��}�l�=уаى�k�|�z{P/Ρ^��~���`>6w��{|�$|r�2����~��o!e+H�
��oű�~ +l��o �Vo��^�xo;,o�q+�e b���LU����Q<��c�%-\w�xr�A�9!bC�W -�A_�bXV�%҉4�߰�]C�R���.�@��y.�����#� d�Zu}x��"t�`=q�$�AeW�wI�A�!|
��5YtHZ�B��!�L��uؖ��Y@O�@W���UK�2�F��4��@�Zb݁�j9ܥp��3UN�&�Oa�(ل�k��-�XrP��85>E��Մ�P�B-�r�N�u�Y��d%�JΝ�fg.�_�n�~���$ �<���gC�/֫��	l�+ւ��qh�n��XRch��`$q:9/& u`B�d[�(�: ��U�{�����+���DyFSg:T-��>)ާ͢�}��G�������"�T.}�R	�0n��lr�RaP��.��g�?�����ѓ��رC(��xX�P��d��HX,SG*i�q�H$b�pM��Y���>h8M>\�� iDd�Z���6�j��-/��x'����+��8
);j�hP�x��GxPuq��mJv���[qx�^<q߃��@G7_Awg7�����v⵷ފ:Q��U��.�C��ނD�>��;3A"l�n2�"��:D!lY�����}D��P��2<�r�n�0�S���CD��^�²�N��o�m��F�9BU��.ۈ#�6���,>��;؊����^p)��o�Ƭ����<7�3��,����ut� A��N[V.���V��h�zQ�26=+���(���Wŗ��[�S=p���ǋV"�^g���}�k!��/Ë/ٌP���f�cE+���ny�8<2�E}��"���{���F�2��X�iֽ�u�{�9w��ܨ(Ξ� ���P���n����^r=v8�\ͅ��C=��Z)t�,�m��Z� d��������7�G@�@��iτ�,�=�b�O4C_�pt*�"���S(�1T*�B)��5x���B�)N����j�A��^ɸ��=1\�q�����`�@7�:�`�:ئ�Ta��N1��;;�"��l W.cߡ�8xd㓳����Smhv����\պ��GǑ�)A1S����dOJ�:����ڴ؆U1#a:Y۲C��TD���t.�e�.;#ݱ����[���D�iQ�^]Z���Dw��u.�iŚiT��p<�hѧ�'�sIθ\���"�2�i���_��4�}-�؊�?*g���xDX.C!���E�������n%�7��f���oE~�rӧ�ъ�j�*�'�'�xh �)��'b[�=2���L�� I����5�@_�tu��sS��
���mk�n ���R��~/�9�A�V�ȡ�0��Z����1;v1O�tto���LzȦ��Ǔ�+�g3���o��T3�B��l� J%��I-�AԾ 
Q�bY(��R�5�L���"5Fgt<�4M`��s�Zt,�T[ �(�|����h\>��8���r��u7��͋�\U�����+)��&���W3�;�� ���F�o���fn]���=�ڭ(�g��po�rxvV8"�O~�/�v"�����0q����[�'Xaȉ���1!�8��>�I�M�j	4\E�P�ʖ��	ˀ����*6-��'>��`���(�����ſ���ԧ��D:���`��N�����c߃�8�\��x��\߾ǟsr��c"?}��!pP�n`.7�G�1w�\��fS�B3#э@�!��A<�乕��p�涾�]@�G����������#px���-P�;�H�8|j��W;ǦQ�l�(	�'2��.��Uǣ|߅I�d��t��� l�vi?6.�A_���,�twc��~���M��琈=�'�!fgsݽ=HgS��j�Zh�4��2��88r������8��ļI�]�s�JNOP�4a�,J'���Њ���_J���r�4�2a�6��% B�Mv@Z d�e���T�KQ�ԛ��!iu�'I�J�0��^O�(��\�uT8��S䥶�kͨP��M�)I��G��������2�zFT�!L ���I?� �>��^`�
��
�,��m�nK;�U�y@(ۡ3���{9�j����@nvcGGP*�q���\�l:�]�u�A@"Ɩ�4�3*w9ئXӐNhv��������1m��(���P��
��&1�V�>���K����aA��hN�0{�$N�=���V�PC��"$x�g2��0l���f .��D��T���9�ƨ���;_H��ߕ&���Q�GdU�{w��7|�e�k|HK!g� ����24(A�^����0.Z���17�-K���'fĺ���-��=)n���B��:�X�n�P7>�G��NE��+���S9�&����%|�h�{��6ztZ����8�0�_�U�{B�Լ�ݸ�K��|�`�8f��Lʹ�ڗ�M��'���� �\��?�N�ħ��K<��H$c0�
.X݇[_z)F��qH�/Ɔ����-/j��ϹSQ� �NY*n���#]�\�#܇Be^|!�������dv�0a�RHe��<LXIl�zy{|���@{�~#�>y~����g� !, ��l�M�����(14|MǕE1K-4���nf�h��8�
,��V���+����u��ò�¦�jq��)<��14YD,8��2!FG�A�Uض�2��z�ѿhݽ�X:�H������>�����؉~̕��]��(V=��uv̢b�����M��@T�1�
X��	�-�@�r%)V� �2ͩu	Y���*�鰟�HzҀD�[������:)��R�E+�p^�Noj�p"���9���"|�g�(^�����`G_�}0������a�2-P�QL��
�0��E��+C&� i)8u�R	��R�B�N����������0�"�Q��`::���`
Q�� M�P蚺����b�#;�3_��TO�����c(���ؽ=p�t�i4&�hN͡rb
N����w�v��iJ��P��Q(V8�`	�"I��>h$�w��1X�nv�h\��MF���������qC�����!�"�9b���m9��|��m3 ^餆m��q����uh��P�.�v�����,v9�'��3Չ�B�;V<lY>��|���^U941!˄���q��ٿ����f��� jkp��H����q�����׮�'����q@�!����J�ͦN��]Ӱa�
̠�*�ǿ�,�F�`y_�r�#���?��P���R�5�-������Ǡ�.�ן��ۮ@�K~��H�'7�: ��cP�:B���ʖ��#�>�S�N���/G�(895���"�ꅯXl�Lu�8�� �?y0�o^�@����>��?w�s��7T��6N櫸�a<��8*"�+b��ET��U�A�導�^CP��a	\}�Rt�u��N���Va�N�ޅ��G�����&���F�2�%��4M�"���n�#O)ܪ�D*�NH��/�֫�Ʊ##x�}���ǐH/�#l���@5�(;
v�>7Р1��0�B�taЌ�rZ5v�´E�
�lQ�Z �(S- � |Px�U���tćj	�)h��2-;��:T�J#+E֖Q #�aӯ�ȠD��rD����� ��5�W�kZ�&�f_z&��U�a!�9kZy��
Pk.	dhe=` "ER�"�&�,��[��Z���{��{����q�l�ߥU����Wb��Uضe=t���SH�H���n6���u�ɉC�2G�#��&Q�4��,S�r���y��hZ=�LM~ �hh���4.Jz�]S����G��O"�ӏD"	-Աnx&��/�`58�*z�A4iz���!�T�5����&��>��γ&$h�a$b�(ۆ��8�` !� �E�mn��Ѷ�.$
\��I>�Dk\���;�g4��� N:Z-�I�!����=��/�{~�:�ZѬ"�X�WF�B|�K���|3�*�=�b���F�Ī�.|�C���letnNи�B��'��s��ᝨ۝�̸4$ �8�V�Ms�nhQ/�Z]r1�{�q4�u�v�q\�ng߅f�f1�����!��᯾�1��T���ˆ�����}���(�{1���^�Wm]�{@G:�����#���=���<���	��1eVR�4����݅�cX�~-�WЭ,B5�X�v,	+F�*m��=��2�=���O�_p��o{n���CG�\��b[q�%02������'Q�, �D+�D� �6-&k����BiV@���K:q�,�_ه+6�ǒ��������$r$&���E����+�$H%�?=O�k�\FgO7f�\M���׽k6l��������׿�L��jU�D��`���4i�ބ�J�)3���Ȣ4Zu�B�!� 1HNYRu�rǢ�#��]zRSY#Mr���	c��D��rMh)�W�urA��R\E�,>f D%\K��}Hq��p9�BU'�(Z�:Fo�����.ԙ����z�h�5Bz�VQ,W�e�K�m���"P*˕���,�K� -kف�^���/Ɓ}�0r���S�J���.�Fٔŭb�ʥ��r��L:	۶H����N|�>���?{��g9+�yQQT�������#������$��/�Ƀ#��F�|�uN.�;9�d�-�[��F�t7r35���A��	���d'B͒��� �"�3M4�v,�KD)oQ�������]�B�P��$�c[b]S���|Õ��m/'�8��,�@�<�� ����ރ���	�]j��X<	�i�²�����q͒�rt������Q�u|�ο��/Շ@���tnن��M�*��`ڨU��h$R�H|�0U��C�z&:o�|���pa99 7l�UF&��ʁ>e�X^���?��l�+#m:x���Ǻ�N�{=�),^>�\v��sω Q�B����6�c�ÑC�e҈Yȕ��DB-�d�f<	M7a.<��v��\tگi��3�@��iO��,�{�r���# D�! �ОQ<udE�4 �Lp�@��%|�P�N�?�㊍k�fQ��w(�c�]?�c�� ���u�lE7���"���r�eNX&S��F��g)T�Q�Lt��`�:
�9ԛ�]ݸ�ʫ��7�?�ۯ��2=è�6���c�/2��J�*���h^$� :ѱt(动P�'u8a:�l��g�j͙$�V(�څ���� �!
ы�H�� ���*��Q�}��;.�{�u�BA;��(`��1��$��na��1��uL��9�Pv��L�&�H�'iIF����D�LL���iTΌ�m�R�R�b(2e[1t�t���֨CM�zM l"#kV_��,��Z���z��`�m��:�?���#�C���avz��%hL>�h�۔/��S��a-7i���MH�Qs��HE���=�)0��M �<He����|�B&݉F�At3�lb�hv�ǗD���fi*wv�D�f!���ZUv&4�6�F��j2 iN�,���\�"���]���Y>�k�ht
i�������u@B���x^}�y����]��(Vz,�c!� wyhj��@1�a���S)�J�C= *.p���?޾a���vÄ_orb=���u"�N��z<ςjV2����gMֳ0�    IDAT�݄�Y j,o_��G𒋆�ç�Ś�C���������NBt&|����X��;�0� +�\�M�\�os���:wT��'�Bb���9��9����#ӑA�(0bij��F"M�tӂiX������ۮ �#��@��������<���hpҵ� !_���T�8�]c�(x6JM�LP�Õ����N�E曖f��Sǋ/^��.[��}�oq��(�	*j�
i.	���F>�̑�)�T��&�T�[\�LM	��j�2,����"|χ>�f�����_���E�ҍȕC�J�s��="�B5F<��u��B.T�񠒎:�ݶ8�Qv4���⎻�(0�:DC# B�J������6�,mw�T檟�P���:��q���S��.�8�V� ���S�Z����@O�C,�d�%�%]�N�9Y]�d
�� �/V�и��r�U� ~8�
\4K9$5��T�T(XR����Va����t�JQvHt:%{���a(I����!@I��Q  B�/.RC��y69��5'F��{	\P�qhu�hZ`����j�8~�5>Vt�i�	����T��C��J7y.'@�T��-$@#��!)C"��"� ["���!}���4���� �n��oe�hc�h�	���)��sGJ��b���h�C��B e����L�OH
O�8�Y����7��GF��/��u�bC��@�|�"�l|&-=q�����i8��V��\�}e���9�3
�w	��
Q�1�P#�kv�c��s'��f�Z�|��w����Ǎ(`��	 +h����ן�c\�!�<qR�[�D�5�{��=v��/�c�p'����3�Z��"��z9��m��s�T�������D��l�) 2��ɱ�x��'�L��	�Hv Fn(�W�x�j� 9�m;�v��,�{�+����+��W<{F`ϑQ�P7�v@A���T��G��Ď�I��,:�)ZQ
w"�F�IK;��qÅ�q����o���i��t�-v�#@����*1v
C��(T��*)-�j99��O����C��*Y�jl�[���b�N�P�q�Wb�歜��o��=u݋�b�(Pv��."_�≈�� �I���?a�`�1��svo��TR�b~)�Vn#�B���
h�LPџ��@�R�Tkv=�bYdS���-}>Y[&�<6LK�dy���D+�D��S�M�0*�Ɂ�4���ND�3,(�FFԊz�3<�T
!�`T��TV�pwGSM.<y軨�Ba�����iL`C�R@ҰPɕ�?{�&WY��ߧ�3}��f�酐�TE�4xA_Tl*PADDTT�����i������d7���˩�w�~g6��}����G�2���kv�眙����x ��t��
��I�M���w��#fy\7`B�2��٬����X�?�AdU�J����!�A��;�L;���lN��d�g�Z��Œ4�7��a B�F�a�2]њP��E��d�o�@9W59�+,�)���2"tM��L.å��C�����I�ՅO�H4����� ៲f�����j@� c�x�?���;a�"��A�,�WE<bq�|?
�2[ې/V�ʈ@���@	�t�,;KDt�� ߿�3u+�%V�#R�e|�����g�Bj�@՗x�<�����A�����'���j�[�r9#]S^4�!�DQ�H0i���n��:b���1k\��u�,>�ٯbǮ(��q�&6jX1����hJF0{�Rtȑ�w�%B���$����"G��H阮d��w�����tK|Y�MA��(:��6D�4$E��H&��3kn}�z�|�׏�u��7�����߻������Ug? �;Zkv�M=r4�2\R�m���b&��0��Űpbo?xN>j.���|�hm$Ͱ�����S��*�c�5@7�H��X{K���֌�]f9��Ij54<���>���ސ�T�|�eT��J�
��%K�A�,C�����-�C�3Q�,d�F�
����w2j���v�ŝ��L-3�cD#�i�$օ����1_Vxg�]ץ��0�*�4l�,/cOE�ʅw��zȤ�V��x<�S��d��¡4�ǿrO���&��chh&��Xht��L��X!�=5��K=4�k:��$#����͡��W4�SK�K�LUF); M�Q�e���Qʻ��%X&��W��>V2��T�sD*��c�>�h�%:���ZB�X�j:'f��\�W�%�x�ÝbdhG=`s5�%�:v��^������e��/4u�����qYR'�DȈ��aXɗQ�׎n0zbC�m�#QWI�H��cϮ���ˣ*�� �g��8�$��Vx���B���h�&�72�@�����.V�X�W ��s� ��+�@(�Lf�F�#����0�G�?*E�k���PY���C!3�� H��!��h�ȼII�2�GW���.���! I5#o;����$&�6#��b��|��`��P!��s5��%�������%��Ě��~�7a`o=h����*>|�g����y�5��bbɴD�>����/���G"�Yg@��et��V��̑�},MC2Ş��������71(�Y�)��D+R�氈@�0�xa�	����]�7�
����Տ�����[��R�a@�bc_���/n�(^ U�mhX4�RaX$�avG�]1���c���{�zD,�����3Р� C�����ҁ%KW �lyf����{�g�*�Қ�ط�� ᢣ%�j1ˑ�--�ܰMއo;
3.�3Ͼ�;�}�ֈ�"PpM�:زc$=��d@%�@��@L G���)7�P��4)�L����¡V7,�bVH�DR.bE���}����Dz���dMf��r�� $g�r?ng�<�ր@("9I�'d�$�kQ<�?�F�
_(�5��I����Ѻ
H�C�;fc�<J@80}��18��g#7:�^�H�L�� �TJY3Ls�3z>¦u	�n1�A��J����%�ƌ�<�筙�k5���])�M�=A�Rl�qA��Q��ZbK��Xb9���B��������$u�T�ܑD� 	�������r���{B�sd�7H#*1@*�3ᮾ�m�S�9sVC �h�MgG�-I��`��j=/�������@(��9����FLԫ�
��|�e@%�;EE�T`���4WDiZ|<2�Bj�*)�]�i̚��ȗ��.(.0b��u?�}O<׊!�%�t>|�I�hL#;4�{������>b�f*�G��%-<���w��}X�)3 �%^i߹�Kx��3���ٍ���_�~�r9�$�hk�1{B
'7 b*f�[����#9��w��}K���E��Y�Y.����زvV�|
��p$Z����DPuU �\I��!���%\ҷ�
�?����~���
�� 3@̿�+���@yM��?We �̆n�W5�z��ó+��
7��	W^|>�l����;���8E��1�u���0#�0��/E���+۳Vl��"^\�W��,���ZF<�j��n,Y�ǿ�|��K��V3����^�©.�V
�j'����L0 �A�h�Wth4$�dȳ�V�0��M~�K��Ė�fu��i�<��z��@��*4��/�2x8��ɕȔ_,�C�!�-�c1�Ɍ�\QR�؅Q�����b��X����ƨY���v%��Z��\N�<0��G��#HR��C�d����ԉ0m�t��f=~�[�}g?GS�S�Є@CS�pXVC�9wɫ:"��������k��v�ig��K�jQc�l��FZR�̒q�ַ�?֏�R��0��2��Z���֐$Vc���E���tH�p��Ob�or}���0$���b�=�d2')�>"&��Ę�"L(q�D"P�4l�P��-N�
B5�+z��x�7���)�N!�[X"I �������1��t�9�."$����&B!����l�&��ڡ'H�9*ؒ&�Dq�e��;&��]�A�9��q��57��<�
�FŞ%�x�7�xV+`sc!j~h[A<�������D8�"tC/13��Q�1��(֛�:�MTp��K������}�ٛA[{$?�ִ��:�F*��k.,>s��@tґ������߳�/�.!�H©�іNB�$<��#�ֵ��f�P!Ś�����m�H$���@2j��[~p]���~��W_��_���S������V`KW�����#ډ��o���Woų�`�� �Pɚ�vЂ*�Rs����Ѫfq�onBז��hi�iEY�Cs'P0o�aX�h�����B�q�oA�4���I�B�fU��x"�Ï~'^xy;�za3��ր���U/��Q��J�1 �K������!�y�)�q �T���TL����%P�a�TD4�nF���G3X�aJJ����9��SwuPҖQ����s���ƍ1�?=���̊d:4����5u�������C6̛��-��_��s�d���G�X��{8�Mi��	㘃dI�r�����IuE�ʤP��?]!��_��W~�gqÏoGѮ9�iM�q�!K��10A�Q{,�b�KC�k%+a�0�*�a<-1�78�"��oej�=4�����O�8z��$%>j����~s=���{E��.I�ؓDq�c�(ò�# ?<�ܨ����̎�d2�Sx �\�\����J:c�p�Tu���*�1�V�S�G��1��ߛ�k�^gD'��!�X��*|�Z9&�Uc���+��^�~�J�i�B�>�P�H �	%\[bǨ��Ǵ�����p�İ�|�p�R��Q|�_�gV�La���^�m̝��3\w�5Sӊ�°߽���c+![	x$�P�%ݹ���O��%��Lhm���� ��a!�A��hB~�\Dgk	���SӘ��B�s�=w>�/9�i��?μ�� ���"?�/�kr�,%�����7/��Ɏ ��[�!E�p�8����6!�n�1G�����Vp�aG����t����_��7Ͽt��/�z_��==�oh UڭUI���g_O�ކ�]��+�̀T������Q�y������x��?A�i�n�-(�Wc ��q|��CM��eV���y�O7���n�r�ޱ�͍(�r0L2��H��q��e�����p�4F+:���c0��c���hל|�d���䯠Xx�]�$0��G��.��EsgA�hs_@3$6��oR�._��[��ß�
�^ڍj��Wh�w���}0$}q�hN8���3��-�z ����Z܀�Q飊|��ր@�&bA�����R�w���҉|���7�ѿ>���!�N��g��s�X����(,]�F�*���9�!*u����LkMJ��v�g�KI[�2���������|�[(x
d<��"|	<H��&y��z�ՠ]�<��%�=�潡!����e�	�r�9蘨���:5��� y~jw1�y��8�\��	�n<I�Pα���D���ꔺea�Z��B�|$��0��"�ɓ��.�XW���4�����9J��xw_���%��..�NZ�:0�<�,,����1`�#aQ�+?a
��]�1�:i�_"qr{����48�M7ُC�I�趢�t����-8�l,��S�1�=��}�B3>.��վ�l�j�ڟ݆�<�"�$��U|�����L	sZc���~aD����ʉ|�\h�&�U
Hc�`��ؐ|����O-�Ue�c�Q>W�aD�@��*�d��&b����1��FP���y����a�ςd�%�� 3�I�F���P)�8�TȠ��	^����+���Xz7ZQ�j�Ԉ'��M��pԑG���!�;�΀���
��+P�`�gW��{o�xn����Ѡ�E����mއ��*^���hp�w�/C�3�բ�������[��aP�%	hV
t�Y�K�<�5}������ٹ}�](e���eʈX*�GG��>�o���ϼ�Ɏ)q4����'�,I�d�w�����`Ңk:�D����Yk|waQ�Da�~�b���Br��$�!�&0�I����ȗm�Zb����×��C(V�+pO����C#�����O��s?|�N|��������4�l��:e��Gc)TK�O��u������\������
���>�6��,_p���O`B��7 SS3�d/��D��UY�HlƦ(`�zOk�H�Ox���M�v߼�	�����m��v�͐$���='dXE��v�G��P*�I[���;1#���>|�=6\��C��NF��P>&YJG˯K@B�9
����B��X�[��`E#��ε�@9��V�� 6bd�;Zdbtj�/��
:n����r�E,aI��$Sj�	t�9��E`!d6(B����gI��#�''���a	�E1�>��r:EcyI�gP��]aPP�؈��\�� Yy6*% �I2���A��cE��T]LiM��o~�����r���KȻ.�������0n���h�|��Oᤙ	is����̆}�"ڒ�U7܎;����Q�kH^(0#+}�G��E*�f�]��uM�M^)�D.�(c|{鸄��,/�V�1s�T̞�M�C��|M?s���{���(������B�Lmm��ݍ{ﾋYk+�Ɉ�#M��W[�/�c�4q�
�(������^F�F^����W�X���k����xS�����D�R�OFUG�g_/o�pE�8^[�Q���Q�(��M8��X0��3�	���2�ԫAO�A6RH�[���c�:e�k���]#�{�c���=��e ��۩����~��x��������lC>�`�h`Î�����Р� �bk�lKs9y�u��}�E����&u�y���Qlpٱ��+���Vq퍷�����l�i��Uej%�@�/����W~�z�L饾�X���_�%�}�i����VC��2\h�Ь(�d�V�>��w�S罏�⛚̢\��_�U�|�5��]�/<��sU���f_:��|�
|LjMI��K�J��p!���d�zfP��[�u��,��brt.������\n�!3�� ��%���@d,:6d��cL@M����X�Kf�����VrQ���~�@e�Eד@�F���}K��E%���Jf�:ڐH��e[�R�q�ZE������D?�ɩ��)�
`��Ñ�v>-�����X���� �_���;0^yk��W�F����(1j��*T-��P���Ӻ��|�R˗,������X�~t3
E�1S��PM.�y0H�������S�)���õ�]��Ƨ�J�<)�����u?�^�"�t\�bhO7N|�;���O���*��X�Gl��h��v�+o@�Ɉ33����t��]��3z+�U�23U,�b�Mb Bó��hm��9��#^�ѳ#0�ALj�y��e�"H�ٯ�g��þo�JAl��1�E�RBDW�И�����o+��i�`��!�	���z@����3�5!V,[�X�"��8d���ھ�o����[W�����.��_�+���kE�P�P��H���VoG�3�aoY��pf�\BgB������w��~R��-	��9��xFs����#���g�W�D~d/J�A�ܲ=��Cx%H��q��'0e�l,?���M���k6"�1C%}#6���@²9����0�1T�'@2�dŁ칠 ]�R@cL��]��[,�����͗+xl����ۻw#[r�l�ʞ	�M�d�&F���&Ar���?���u4)�潣�J����{?�y�y\��&<ڕ��L�P���Uq�7.Ƭ�- �XԒ�~�r���%W�$��D"b 3�;��9�݈Y/�lq_�����hH��eIt�~n�_�w�B����c?�+�JF�@C4݈R�M��P�yf�U���c���`���x�톽��4�������Z�0˶Xo��%AЎ�J�����𪈥b��^.f1s�\�q��    IDATt���<q�;L�����s�B�cP#T�9ݠ!?���$Lˢ�Xp��h*�r��� �D�J�Ymg�yI�T�=Ecѻjƾ��	��j�l��u�I���E�,�S�������Y������{T��݆�>��G*�d�d#��J(OS�>;��M��P�u�4Eu4G|�k���3���т�\�ja S·��/mۃ��`��i
��0Z4���,����gXV#.��xt�DRm�
#�R��Z�����4*Τ�zf��Q��&y
����� �2�up#D��,Z�)�V��}�؅�"?: �.8�g����;U�x�O�p�t,ـD�D=�m��р�Ҁ?��z��p��C`�%�t�@^�_��czì@��a.U�@�+�q�6��������d*y|-2~�� }�F�0D3[5��t\p���+�B�%����hP����p�>��)N+������Y�r�x��`�E�/q��$����S���������@o�_kÖ]9��)��ȯH[$�Wչ[�Z �8�C��LѠ4X�b��rv���̟����K;�Ҏ�+�|��/����!�HsA�_��Ѯ3�*\�� �'ۏ�}�}��٧�؏�}âd{�7�b�p	=�<���<�4�R\,��ِ���oK�O�[�"�Lᱧ���_�A�EOF�$)N��s�  h�.�r��2�p�M8bBRڰwD��I����?�#e�T��!0t�6It�,�S�5�G��<H��h,��+4$.��X��2Ƣg�:�	�YGUcD�K6��w�����6y��Z|l�Bt�	4qY#w���ځS�
>w����'!3RA&oÌ�`F��~!�re|%J�2��¥5���+���(��
�1�K$cL@�g�~������2ᚌ����bn(~�$d��='�+|VQ�~G5�{����@�η/�Nz�l�@97ʩf�u�ؽw�� z�Y��]�O���Cz'�j��s������w�2%��������3��Ew�I-M��;��w~t+�ߴ���#|�A%�<�+.� G-���ZS��g����Kߺ���VC;F�E�F@�2N�"��*��h��g ��J��MA	}
t�b�=�L�ɍ޿�v�&�3g��A�Gۜ�Կ��7�)B%�˫�T* ��#���o/��.���4R-� ��W�hD6���{����N�d1�riC��ŗr�5޴+P�`z�^����3+���-"W�s�,�=_�p�ţ[����>[A�p�W��`ф8NX>�6?����S0���#9=��3���s�v@�g=/�J~Q���C�
t%@�ZF,�B��N9�#��7�_�}/�Zՠ	#e�2Ȕ|N1
B��%(z$� �LƬ̪�A_��U�� i7^�-,gJ�sbAKRjXq��T$��:=��aX�'	��%���i�ra�6t�����u��!
9LnII�{��OaRR���8x��h�<ùljHOD�{�ӷ�ϟ���΁��ݚ��w�_�e��j�d�*�S�(�˵s@�"O����!��{~r�e���	������hI�]�Sq�}A�m
�n �&?�Ʉ��,��gr\���xD�Z.4&�Iyh�j�& �껃#x����әjŁ�ϯz`�{��Ɗ���%(�iyd~���DRQ�G�!j)8z���������1�%�z�H�~�Bt��C���\6L�b֣V(��	M�c刉����^|�"5��̪5�83$�� ���V��)`�ڌ�@�<N �����"��H2�G����`��CT���݉�/�b����"O�ܿpw��]�|��X��y[B�%D�������&|Iŧ@\u��0!mA�Lmn��[�wX\���a�K[!�&�ݰS�އ��:���s0R�$MiW�>1��]��[���m��ɗ0X��X	��l��@d���)���K�9�@��!�h�@@S}$-S�޷�zi7���'⠃�@����?�9����l�A�w��� ��c�����SO��T��#�4�Մ*b��)�-������OĲs!��D��t����;.f�5�+P�).c�$^��޽Ke�Qtxd�T��v`׈�~W�`��-C�a��4N;z�7+x��[W��Q���C�;	��>퀽�r�]©d�F3$����#�#�5u�9,)��X�x�t+n��=�8RF���)`(g�ٙ9be	�i�Ħ]W2S� I-��0M�J�h3&4��/� U�-na��A���S�Z!�ƒ�`��K��@���`��K/�4K�sbzK��k�HE�+Yx����&�s�Ų`�]�MW|��䦊�Z����}N|��l6�V�|{h���E4��[�8a���+����o���Һ�Y�'��˯�=<���Y(Q����R(�"� *=�.�D���Wv�k~��MF�ֺMj���xʪ��W�p�	a�Rk>�� 9���xp��$��rA��}-�t�@vKx��+p�����	���gȄf5 � �����O|��;mjE��龨�b%�@(ˣ�G1as�`�/�%��xyc~�����3�(18������@�����W���Ҷ�Q��qk;�<c�@�$s�#݋*ES�HN	7��,��T|���D4jA�����˧~���!�ؽo�b�A���[C=��=��_|,^1�Ţ���>p��~�'�PI�C�-������>��]��TT����;���~�W���Ӹ��ϡ,T�$#�T4L4�&$n�vIGF��$F�1���eiPd���Θ�c�%�na8y�koŬ��1y���)�3���=��S�!*�A"�^��JĐ�ư����� Ex��t�L�Z#\%��gbǨ��x
>�CX:� ��������@^��s��W���y�_���W`���D�T�Q�Q�o��g7�¦��r�j���L?�C&&p�Q�1;-�陇�d ��f��<�#�s�}��['�jɈ�{��RX��.b�$�n����>o~}���3RAΎ#0;���Qd*@hG;��~�I� ���\.��CQ���|��)X��{~u�$�-��^�8�B��N���3;��]��l��%�i�I��]�r��7)թ�)`c�{�-*4��o|�_މ��#�pU��P��a�E�y���l0��dRҐ~�����?�-���F9%�vڞ&�o@��t^.t?���]�{Z���H�kWߌ�X[���D).���*?�;A^��o��"�7�X����?�Ka��+?� :�|�5ǘߤ懠1���ax�S�	�IIn.R�8H�wȂ���/ � ��,MB�PD��=e\~�MX�~3��F���'nIPe=�a�2B����W?s�>�8�f6Ƥ����?�iT�*�	��Q�.��(&�� r����y�M\�J�jL7��N����3��*7$X��s�� �s�r,n������,��;a�⦜'�سU` _ş~>� 2�<�H,좗��ٷ1gZ'�q�g����,��eS�ҥ��C��У����&0�,���qh�*m)8⠸.�Έ�Mi~��{sb���tǳ}�/}EO�n�f��H@����J������HQBy��8ڸ)C�ec�t3� ��Ǹ�f��`�Zr��[ۈNŭ�+��K�\��RG�-�$��гk'��	X)$g �X��el���U�㼏���gO��B�T�lQ��~��^_��+p@��:�W���/m�(��2*�זC �q7�t���Q��FgJ�s���٭���ѳn%T��;�E�Zi|����j�u@�g�ݫI��1+}={���e�"fC�Y�t� �w�uzG�z;
~]�t�A@à���dR�2eP�*��rJ�+C��k;���W\���뱴C���$ �8Z�7�+NX���2���]�8u�/eq�����ދ�A�@>r�'�$5�+U,lm�n��j��ވQ;@�m
�by�,���_~�����*f4ǥ;��(>��+Q����Xb�"1�2�0�Pu������'$��}ya&�8�o��m=��䨶�o��(��$k4��~����Q!��EH�C���R�����<�`�7G"�F�{��c�k@�e�Ȼ�J&d5�B)AK,�����Ƅ�F\u�Ř��(P-���܄m]=x�ѿ�/O>�����2~*���U`',V$~�1�Pp�� ���{�Řܨ�8�M:����-�+��wn�y9�F ��Ȃ�N�
Y��-�(�M��^a�!�
��� 5�:���L(]��xD��8x�4�|1��>r�Ri�HQ�J%��]#���1XQ�_���X��J��1�!��E̢�����P�7�a��I�$�(1-.I[�l!�.4���=LM��^��p|z2��\��]�}���3�d`AV�S�r�C!	&T�%��g56H������B�@�ZcvH��(!�8HF4�����������z����ov!Y�c¯B�%�+%��ql\��>�4�1j2
9Ҁ�H#�ZQ�x�{��z��T�3NƜ���(�"�:|�[v]_�׼~lo���y�ש~���X�a���ʎۑP��G�ۀu�#�Hq� ��A��%�m�8��ވvi{�=����s��I�r�0���[���N�w�P�"t�ņ5��c�f8�"�4�َ�xc#�O��F���O�@1H`kO]��aǟ�M��0#,Op���q�Qm�e��#�	�Tw��{8bJ\�QB� 3��ƺx�:$H6Dq����q�D(I�)���|�]Kq����9NWw��>�:h�|�Ri�p^�iJH�����7�yf-r"�x�j���p�w���s&B*���H7����������P����n�I3!��@ ;P���z�}r\ڙqE������s��L����iǙ G��-�cE�w�82�A�˯�	c�bN���(��k~��p<.K����>��x8w	��N�G�Cx�+}\4ȏ����RJR��ьݛ^���};����(���  (������\w��8���c2ʾJ!�
�|)Ϭ�H��%FX�@S|X^�$.����u��A"�Ƣ�ӥ5�U�سk���^������$˓�yt�Ċ�Li��Ѣi>v�_�q�z�!��flgE��kK}%��(F�� bLlI�9ia�����]�i0'�^��$2����cJK���sX��M��+G	 D̸��?G�P��a�O��:&7� ���@ALn�K[�	z�i�ii̸�u0'���'_؀�n�5F2��fh��1��7;R	�5�L^����$�>��(Κ���H�Et�l5Р�H�2����!G����x�7C�����KG�����<��@��LɃ�W�E�����-��f`�&�Tf�Y�"x)�ź���ڟ���8��0r;�jR��#;p�"��	�T_�7�
�������_�m;���|�n�(]8r�<�<6��c0�P�:��E�F��3�q��&�W3ص�)�d�"C�,��&�p��PR��xt�f7�Σ{�FlX��u�4(S�e��rS�<��*dф��Fw_�=�<Xs��	@7I%�D��4�
�P�D��7���\��M��5�	5�`�!��7 ��,n��?d@��N����u\t�ix���!����Ӄ�}�+�;1�u��1-"I[F��Ƅ�\_N�r���㾕��[`���n���8b�t؅�h����r��'t]��rf|j*7�I.t7��]���p�D�2M�w�X�n�d3�gS0� �!�X.j��1=U-����N� a�,�b!�!0��o�u���΃���?N�Vu^j�=8��Q�|m����s!���S���U��t���a����݊s>z:>u�Y��2��C��X�f��a<��s �mlC�P�r�<��.>����p�:II80hUs(�x��m���;��܈��mҦ}�B�&���~����@2!$�{jH�')��S�@�kQ����	�*ޣ�
=($S�0=ʣ{�X���Tx� ;�/��O���~��
�h��U	�S����0t�]�@����7�="��X~a2���~:Ύ�}BeO���E
�Tn`��Fi�ތPS�^'�F���n�����{�w �h�1.k$`(��<�'9��J��"�ot��# BkC����/���7�� M���8�B���w��sF�ǽ�z+��m�8:Ϧ�M˄��(��?~�H?���Y�%`65�,E��,E�s��5��b�h�)��g���C+ea_��>C��_��g|��@���������V`��-bpt�S�IG��#k�qt�����VQ��v͖���5�9��)b�KO!.�P�Y���V������v��g�����!�y���]�7cˆu(�BDSu6��7�b��-,K���I)t��g�w�i�����H:ſG����j�[gF�Z�I,�U,�=����ej1�@�Z���B�y�%	?�$q�.��!�f=n��wМ2���d�8���"�Ќw���8��w�R=X��YMi鱮�~�t;��A6����h�TK����$�����3_�Ab�@h�<�҄hpW�QZ���><x˵���{P�t�+o��k7C6bD)���\ʱ� �������@�^���a�,f7�Ν�b���;w������I��,�SD"K���IKtm�<jE}c%�$m�'�@���)�0܃9S[q��b��0����e��2��;���!_�@O�����.b%8�6P,3�a*-2��u��<t�m��)�-T0�9"m��-�N����p�8��s �&���A�iTU�s/�e�$�
Y!�	Z�Ğ�7� H�(>�w)Fׂ_)A�D5T�N^9ǒ���F�|�/Y���f��-��%��
�b�}2�X��j�ݯ]Cbl���6����]#%1�1��-	
R�ŝ���w=��+ð��@y��ʴQ](p��!�|+���A�	1%�K%!����
Й:S:&�X0��<�0̘9���h%��'��4�>������������rLEp�
�v�����v6��o���m�,�y�$xz�*q���xi�0�?r�@�}"�Oj�Q�!��h�[�[������z���[�C�r1����_�;v���~N�R��̠{_�v���m=�SU��B*�Ѩ{X:�G�m��D��>���Bv��j&[p�韀��������m~rP����>���]��2(���6��XlE�ֽ���-�x�4l�E�l������N�bV"�>a��@hܑH�%`�fOn�m7}� ʥ2�D�8����-6�3 ���pX��U00cB3~x��X1N�vU=Aހ/}�<�j��Y� �������<�^47I�^��ܚM�ڳ���7~�RL����cvs��؎Q�/~=y&Khh��|tUxdi p�Ĥ2��uX֦K]CE�Q�r�Exy{/⭝\<HCoX�Wۉ�I���L�<��u��|
B��<'d�j����$����zП0h'}ܸq<��޽;%>E
��M��VP�P��]��I��j�o[6_��98nF��u8/\ہaƑ�e�x��4�C�j��V�n��: ɾ��d�?��L��z�*��Y�1m:E�%̚ځ3N|>{�r�~ya�v�H�1��M�R����ۻV◷���6<JG�=�;�llB�P��c҃ϓ��-��њ�ȡ	�c C����I�x�i�)Sz����C}�����?G��X:' nF��p�JU�.af�)ud��k��)m�RW_?_�)a��摪��`������Qx�
>��iG̓��
����O'=��Nq�5?º�=H�L�n�XB�Փ��.`h0Z �L�{U�� p�`@���kE����0%�R2&6���6�\$�"�Lh�A�g`�E���dXF���)Aa�K±s�*Gv����UDLz*���]x������)�x��f�8v�(Xߝ�ڝ#(�*L3����矊e�
    IDATmq(�Z��: y�\��q�!W�@ސ��~�jv��%z�+�y7U�l�5��z���n�s��M��e���Eӛ�'bAS��BT� p(m%��h�)g��Xǒ�>����0d�(!Uеu3�Q��ۇ\����apxц$\MǞ�z��>�Ԁ_���h�M��0N��t��ƒ&=�,hJw���A��S����q���~�Fl����R)�'�q�4��]
%K� �1��/�$fLj�W-Ê�q�.����EO�V���;��d �D:E�*~u�]������G��|�:a{(z[v�������DUh�U' �@�ե���@�9���M����w�*@��EWa}w?������fh���0̌��4�U�w�-�v��;��Z��r�٨�Ɵ���Om�Ĕ�T.�� ].����I�^%9���F<H����� ����4v�_�\q�1Ү|YLJD���bNg�� K�8	�~'���l��t��zu������u�1  ��Y1��F����z/.���r,�L�m�'*Y��@ڰ�'<��F�߲�m�+�P���D�(Wm6���b���ń�E�1v�3��3��h��4�s��Ze EE��r�x�@ntɄI� ��(�,�'O��;HG�s�М�A��OiMK�����>�QT���p�u?��h�$-U7����&�O�w6�t�
i�pY굢I<������7a��sW�j�Q�d%�G�*lj��\��Hb?H6I�G*zd���ߨ����r�L�פcڤ	�5{Z�/��)(�%4��y�y�{׊Ri������QWO2G�2 CƋO=�u�֠�}<F\��vTe?�=�:_�뺇�iM%��}�'?���ÃhKİp����~�����[_���
��<��+Q?���
l߾]�r(;.����d�����]xj�n\)��.bjk'9�t*ظ�O�P�A��D#ֈS��$R�Q1?�K2����wxE����{�ª��p�Ȉ����`Ɇg���5�o$��}(���fJJ�
Ŋ@5uPSC@j�ДZ��̉@]�����/�!�®�Gb�����jBw�@MC�����I�T��=G/�w/���B5*"�4>v��X�u z��bg|�m8��S�0*K3Y1'���2 .������U_���MŬ�F�L�c�6�/��7�B �qWq0�%t@58	K�G��m���q��=�T�������^�B��e�|4y �1 ���X֫o�0k�DJ�B�j���j�
A2�k;�lV�Il���Ĭ�ᾏW<8ܓ��@ʑY��N��,�C��FJ)���?�'�o�6��9��K�z��ٝ���w�_��-h�4V<��;�ꪥi�Eל�wI�vx�7�Ϗ���8a�Η #ŠT%/$-��5��K>��M&D��Bq�t
�*�%�2n��i�~ןP����^-W�j�Ybe��f̨N��c��J
�j*{^����n.!���\#��h��ZB���f�Ea�@��Y�1f����Z���F�<=,5�9�T<��{�CO?��<+J���]����5}2�;�t�l
�� �|�2l�փx���bX,��ɟ���6zzmj ë�6�r7����\�i�q���H��5����F�ރ��*��oE{�8,Xv4�h�����w~��l��DP�f�(����}S{;�7�=��f�j��e��:�Xj����i�#����}ȊR-�H:7�Ϟ�~���?4�清9���g��Ů��z�o�7���k�kׯ,Ga����:
���<���r��!�+�K�%T|蘅X:I��'�FZ���\x��Y8�����1J���d������|.�S�*49�����U/@�.�@G��"v#��Vr&r6n�Ǔ�T���S��B�9x���\rW�`)%y>b�	e ��.�Q�$,8�dD'Ah&�6�h�J�B&@�,f@�����΃�ڨ��ȕ�s?�Ml�-�JwB7%4�|�3g�%31Է�M萶���W|/��_���Xv�B�Q��	��׊/_q*Z*�DЉ�y8]��! �}�Z��x���=\��bґ�\.���- 5R8�sK\x�ю*k�j�����ZNŻ�^� 0B�jE�/���jC����i7�@��lb?X�6���AR��e��k�|�� {U��e������R��ߛ9nG�~���/���Q"�y�݃_�p"�R�k �c��<)q�z\�M�~�Щ���(F�L�N�(����SO8���Rw�*��`�R�ih��7��'�~�=�Ǜ�/8(;>�azy*��t�1)�O@0�����I
ƚ:2�K>�(�� q@�kG�J1�_�I��E�J)Vץ��}Db�|hAm�̜�s�<G�n狿�/#�HK��Ή���v<��:T��b( � ��t��;hْ8��waɢ�ؼ�]�U�dm��P�`2��ז�9銒���l~�E)��ϓ����49�
��kՄ��7#↋	m	̚C�U@�YƤF�TY�Ǝ)P�Ľ ��E�`X�QȲ@:��#+� �U�y�Y�ڹ��P�$8��d3�������`so^��T34߃����s'4���C�T�li����?�[g� �s��g����ֈ\��C��P����������_�oǐ��$��4��(pļ�{q+���	g-2�J�� '�ǩ�q��k�>C�[BP� bRz���P�	�>�0�mݎ��6�01���V�e��8\���v�屻o�O�qءM-׊a2K�G,��M����>��\^f4�}Q�@s\���~�LMH;��.yX~ԉ�ڧ�R�'��F�q�ڤ&�꾏�[���z&I��ihXdK
���w�}�%����wἏ��/�D8E (�0�5&]��;œ�?�S>p�-[��Xq�Z�_��jd�7�<�Rc2(&� �M.���]���1�2�f��	����T�����M�n��)�@Uh�HI�q���Ƀ`XѰ�0 s��=5z�zB�{,�GB�nH��/4�ݳc^�����wJ�"O��sѮ? �vl=����U���ɺԕ-
T��症�E�^���Ğ�,�F<G�T��k�2=Ӯ���0N��ix'V��!��Tx=U�]�x<��4�.B	n�?��xױ+�h�T�NHҺ=b��Vi}o����&����?�y��� ��Cu����FP�gY�F(
vX�4��u1 ���B�h�2���6�Ǡ)ReA��Ы#y���#��@�$tm)(��]4U�vxK�h�o��/��h
�WCyA�v���?�/�����pI������M?s���K]#6*�I�DEc�-1&�`I4Q��D4QC,I�D�����z��Sg�������Y4�)�W��u���|����~����⤌U*A��F6�լ� 8@ǿ5�3N[�׾�ո{�|�ӟ��R̈��OL�5Ƶ�9��A�?BH,р0����\����|t|Xʀ-�ݓu�`��V���L�<����q˙�x��=��Rk7n�_����*6h�W�Z�"��uS��H
ؿ�.��yb6BR9,���	��kPOҘ*��Ώ�A��Ae
Bocs$�qų��Ӗ��]8��g������K?����
ܯo8K�vi~�+�c�nUi�d"@�t��l�p��c��z	&��	�q��]��	�|���p�0�v���b�������`�i�a���S�Z�bN�:�"Ϻʌ�^\�T��z�B���B��PnF�o�h>g�(�#���?#�S�h��!�C�-��T.#kЍB��YY,�YDێv��v�i�(��c�D>t�&��"�#�WD�Ցi
��b�8��4�U���?�<|�]/C�>�V����Z�����{�`sh7+H��*£����<�)X���M9��x`~^�L[&F�,l+_���?o?fJ:��]���$7�@��o]�~<a�.0w�G�O{)�����(mg��t��H���H�_:��i-V�A��/ڦ����^�ߧn#JQ/�����A�|=a"�S�~�z?���8!��G>��~��Uk ��Ю��M��'�Z\�)k�ydF�
9��7�w��#Xhm��؎\�ݦߣ8�m�sRİ@�<��"���9���.
�*9/"R���l"�
>ڵy�&��,<�I��?ؠ����/��zް���oS��̗1yrn6��<�1)	����!8|��5�fJ���Sz�o��1^���\��׋��?�_��k`�Y�n�vq��q���(<��,��$�۶���I��+��W��\8n�g��Ջm�p�=��羂��0�L����`���Z�\ۂ�ب-L��~V +�/��e#�N��)�e�pC�bA(-3Q�a��T2L\� `O�؀gYƘ�Da����kJ8�8�R�=��+ƑNg�;�x	��i��{aJ��ϊ02��X�<Vi׃��1�xͷ���^�N���<��f���?����8��m8�TہX};*FΌ������i9�f98{������Kﷴ��
,]<��
-}��
�?|H�W+�5%��َ1�p��Y\��f2�=�H:J!h�1�p��q�϶�Cf�����Z��G?�2�y�#���w�gv)�1$��.š�k���G�]��贛X�|f��ht!֛���t	=��j/����8r�*�x@�3(X|&���m"](��a�$� �9!����8u��r��O�E���A��㬋��fς[\�`�;�F�Lې;�$�5\�����;_$�"�~a/z�{p�cN!�EAW���]~)^����gO�N��&�r2���=Sx�ۮD�B������������3/%���f���&֯����؈�z}0
eP敡iAq�ߗE�83	7���BS��nvBQЅ����L,Ezl� �@LAS�!�����IK�ߧ~$��q �u�T��0V��9�?Ϲ�bXa(����Pk�'�Q�~�����☁z����otč�u,���s&��S��9t:!ɗ�
�ܮ|6�se
p��A����v�s��/{��=wv>��X�ʘ
����{���9:6����a
)��[�?�
vj^6�N7�QA�^�����^�x������5�;f�c-zU��P�DX�'QB�ӎ^h�	�6�ay	��7c;�	ے�~��Q�K7�S����b�ܒn��g�ˮz-8�P���g�NyP�/ic�L���&2~�2���\L��K��@%@�V��>� 7$j=��Ng���X�/�,��Nĸo=ت�+
xĹ�7��E�2|�Ɠ����_�y�7gw)���<��٩�Ѩ#��!��"��A�O}�#r�:锄���43;��u��L��>+O:��N"Q1�����O}<�\=�UAtζ���z�/��}b�.���aXڈ��
<:��+eD���h�#�vp��~�� �W��&��V9�Ĺ�L<n�'�מ�G�$#@3�b�ڵ8�c�Y"2|�
��f��_1\�BY�;p�R.�b,��q��Q�(����1<TB�(�[0�<OW�6\$�aTzZQ7�v��3̓E�bח�m�$�S������b
lW�6R�'1<3�|��X���b�?��y����m�}�nS2@d2`;b�T��?���cm�0U��d�����8Zi� =2��b�CE,�8��+�q�?~ �zF��3Ɔ��3�j�ĸ�Ϧj]uÝ��ڷ�QzRھUr9�$6=�����D�	�+_�����r��(.���8Ri��#P�#�?�]�((Oi7,���tH�K�J/��.Z�
\�@�w�X��D6�ğӴ�2����}�+��on/�N��LF�Oj'P)ח��ܔ�p�`�S���v��Q�s�T=�<�u���ѿ�����;�]�F��$	�<���l:��e�R)_��uT*��x�d���/��-[6.t-�K&�K��i��P.�R63	`��mZ�ϝ��P������V���W}擘�/�{����Ms�z�ӯ@��a�)�M��2F��+�K���:J�y�t���Wb�#��Z���C2ZZM�S�}�L��q����;߄K6e�m���'����N�z�?#�����h�%���+.[�{2]j��:đ/ir
��#:dP�@��r��Z�b%f�g0=9%�WLL���ת�&�P�#@�`��sB���矾��2���-yA�l;g�������k �:��C�>Dq�nA�ņuk`�3��:t_�Ʒ0<:�t6�$�AKyh#��*`��:��C�u�Ǘ���!1!�<Q7�♗=g�A:ia4��̍\'���3yi;�+p���<p�Ҟ�O� �\yAS�,�N��r?>8��s��J#``� � f��5� /��"���BT�B�L�[=d�	��E�������#�J����󭫋�U�@���"�$��ub�V��0�F���?݁b�$��N�/`��$�_�P|�t�DaJ�uX��14[�l!3�+K���YG���o�i�a&!�i[V�6�c_���k!.~���F7�У�EM��8I���2��:���g�ʷ��d�0���=���?���Fvl�ZK\�<?�Ab�Y�z��	�z�*�]�3��\{�z��?��COy�����b��q�qlO���j���.^�7v�.�T���<��qh����
 aҵ�ܠ;��0s!l3%�2�ZdN�`ö<�����6�(��]5���ۢY>6�^���t�S�aRt�u'�)���t###R��"�v�6��,���9�vRf����:�p�g�::��X��c�MϨ-�&��s-u���kW���(rV�*��h��EX�5�ɶ��
�M�jMپB�ӈ)����W�z�q����3S�O��+W�����9Պ"��r�|�_��z�%�-�ǠFv��|�?�-�6� �9 � ��c�o�p�����a�Y\���w| N~�J�ץ[�؋�����ZX�k2j�ۂk*�뗕������|$�8�GpͿނ?���"L1]��Э.�M�Ħ�tC��N��,�=8^�nW�u&��d3Y��D�2��b�go;s3�8���F���3mW�$�	��J���`�=�aWa͈��,�b�F���Fyȃq�9�Zm������.E�Q��J����hv�P�lX�F,���6�g�ؒS�ex>RCcX̵mT�iL�u��p����	4�m1����:v���>�Rl]>�,:XQ�a˚_ӿ�}^z��x��� y�ɥ�������Cjn�, �Er[8<_ō{�⇻&Q�Sz�f��	��n���g_��2����"��y?D�Y�������O}�@��y�s|
��#�5�n�	ϵt�byʢ�w,��udH�����}Ǐ��fQ_l���0�q3h	�]��8�k����J�����Z_�*�څX2��i���dj�N�\s�H,��i����|�/ޅ�e�]�u��.z�Ӱz�yht�(�e���,)�^�{�o���Nǟ��+�m�5���*�=\���a��`H��Ai^E�y��cy^����!��1WW+A�ka�r]�^�����b�碧�Vx���M��.l�Vs?���`�E�UE��˞�L�6a������-x��y�&�^�w��.W)	Q���y�t`M�����G<�<�����0��P�u�ֱ�*_�+���{�uu�p�8��PF��cjfN���@�P��H��q����LZ�����Ԗ�{�7�ɇ��X_�`b�lY�T�i���0�	���X ^�`�HI(K�fK�vͧ��NR�����q5[��Ie�/���S��λ�=����:29�����ܢ���-h��O`�]A!k�o36�.!���ȍ�o܄w��0R%�b�?6,Ǒ��1,��:N
��x��]���    IDAT���*D�M�w���5aXh*���y��g���;�Y��3u ��<�{&ep�Hc
�cfxh}1S�U7@�P�kF�]�Z��A�e�d�4��0ڵ<数1R���C뵘 ���c�l�m��k�������q�1��t�B*��Pg�}6V�݈������_�9�o߫�xHEaa����<ڝJ�<\�B�]���l�ò�1��n��O�"����:����A�*��L宏�'j8Y顓�E7l�^]�G1S k&��y���V��
1�KᜭKI�������_�t؇bi��+���~U�W�Ġ5��#�:~�c7�=���[W��J�;m��.b����e(YmD�ǐ�*(��PAFdJZ��kq���b�i��#�f�.]^r,"Z�Lˀg���B� ;��ż�w�OÑ�C�=9)<|�f
�^� 1Qk�)��"��,�=��p��"jM�raP�̦��I%�!~���S��ƶ%�HI��!�2.֑�b���ͯz!^��g��t��N�����?���؍�f����p\��yZ�j0)[v��G�����k����jt�H���W�[w���Ù�$"�D�f��U�|�=�����۪�0�|���eˍ/޴[��-W"H��G:��'1��.A�i�R	RI�\�Q<r�k쨴Tf(�K��2T�Z��?�6����N�+~�֨�l
�{5����b��RN�x�k��K��Um��gv�0��ԥ~�	��"�t��r݈��kr��֍ݫ}�s��rl��t�.����-����v�ޟ�{��r�B�ঘ�J�ޱ����;�Z.� �ayش�7.���Z�v�r�q�6�Д�=S'�[l��<Z7L�QWk��Ʈ�E�,Ne�ik��?�9S�M����^��λw����3\rɣ�o}�Иv�؏�6�7��اplz�!�^�E�
�͖��{�A����w�B�`�����!p4d�%��z;����"��1�2�w�	O�:j�/7i�^~��o�K��.�;
=�t���'r��> [b�w�����u�P�`t�$�.�"t��LM$w{���a����/ٽc'����n�ڢH����ha��X�D�qc�&rv��7�!m�1��1�#�F8��3�v�X�y�}>%�U�T�Y}�Z�h�x�t{��11�^�0�q����'��b��/�@'��XLl�q`��;�ψ[^=�Љ=,�Z.��Sg^�tZ�:�K��$l��"VPʸ�v� �/<������K ��yܖ��״;��U�v��� ǪM ?�L H+4�P����V���۫��Vaۚ
qF���X�*�^�ts�(��`���v�z��L�Lg�ް i��	4_��C��(��hYz�:�Ƀ�t�OĭL�v6:�BWѮT��|�����?2]��89�̢�o�$$�K�a��m�P���=)v�cɄ }%��'=�m]��=\s��O/*y���|����u ��/�ȉY�X�;i�,��D�I��G�����W`�i��VT'���_�C'*0�BCkFA�=AH=��׾���K��:�0���W�/����?߮���!ʍ#���wLXQ(Y�=��.sL���W��ۊn;@���!�y.��n����$�� ��C�Z��F�XԷ���B�"crf�:�^���yx�S��"�PCd`�PΘ�4�Y�]��CY�?�{����N����Z;��Ss�vLO9��j�p֘�5'F��Uk��n��LubŎ��|��y���\^4�L��˅��|�pS�F�-:�RX�s�=G�k�ذ�h�?^Vn��,:Z��^"�����{�ijf^��5�:6��cch�����|���{�މ�������]ظ.�&��=�u߻	W�K_�W^�6t�w����2����/�B;�ti���4R`j��'b'�O�?Z��E��g�
� ��k��Zx��\��k�/��-�� q��tC���нH)���P�8eL����k���叚��dȈ��Iz֬\%��v�N��VK�Z� �0�4�HI�$5$�A�\�b�Na4A�c�Xk�|��aE(�c�2��|<�9/�h��C72�j�}��.O߭f���-9�ؑ�Wo5�]._̉�݉{�랟�Z�N�G�H������'p`���G+b�݌��i�b��i���E���-۞a"�x���cJf�9�W��z�_ӣk�m�V�~�K �~wȖ6�׹��U��{5 ���	ȿ���(�f�n���Dp�I'�"�`�Kp��ql_?��Y����x(��Nh����v��X�b9.xЃ��C�	H�D$N"���%NJa���i�8q�iX�e�`�Y��֍�R�H�54��3�8|���G�0_�+����}p�"�Pb�J�%9��R^�v�pz�� �=p������?ذ�lƎ��*�:�01b��؜J����Ǿ#m���Wb�]�[�VO��!�=�&8s�������pt��S'q���)�q�9qa�8�VF,��@!c�8}�J<���q�c��SK߳V��������Ւ���@�6�"ҤT�`��I���O<WJQ���' FNaL�4�J~���.;��뵣&��&�
��n��=�
	�x�3�'](a��/}�8�UR���:��X��R���Z������z�H�� is�����*����@�����V�Whka'�����uۡy�U�_(��!C)��Y-���h��ey��Çabl�+�{�|`Ae|�l��B��hwC؎#j��p l�Ʈ-e��ӯ_V4�ٳ_�u�fcߑ�j˚��ޅ�:m$g�4��|�*\�����`C�ɏ��{�ðiM	���՟շ��2�,���M�C������w�=�Li�N�P���QJtp� F�H�+�γ[P�NX�����*�������>j�.7���P	��q�?]+6���"H��i�$ȋc'����}C,���3V��AB?�נ����q���>J�����
�9" �t,&܏n����ͳL��/�� a�G��;	�//`�!��2���nM|'~�����3Β�C%��}����NJ�i�r=U�r-i�p]����G6���@u���w݉�o���0���n�B#I���P�0vMNc��j���+�A��Q³riOl�	BÔ���>��ز*+����lX�d���|/��{� ���.��cn߳��}Ć�^``�\�w�:  �f�Bˑb�.�R��C%?V��ʢ���^�s�pt����a���}�!��'9��b��e".�f�"NtAis�b��i����ɿY�Hn��nG���Bd�Qc6'�D� �q�����2�N�������c���� �FÃ��a96V��r�-:{�v+�O�C�'8}]I�;p�Đ��1�`���X�'��x�����'HM��Ǆ�f�"|�V�|��>)������7^	Yd�#�	@�)�����y� �<�t��/�z��������|���G3Ik�.:%�d��&���u6�^�;��5�x������k����2%�!�ɑ����a˿��+�	�dF^RpR3�|�~��l?g3.{�ðn�2)l"��\�r���.6�|�������<�}�FmfZD=�i�5�Px��$�;��b<�����G��ə�bg|��㧓�o�~||����ZU\�Z�V/_!��m P洤��b��u�!���cb!;26*I����
��li�F�����8s�lZ��֎{���Z���Xlu`���q�~t�|���5���t������/~&�`�m��5���z[q��L�m7�� ^��?Fnt5��P+��戇	Q_�JঀmI��K�-a��F�H0���w�	�n76N��W]����7���C#q�D��J��%B�A�[̯ �hX��᧗�E�b�8F�cϿ�t�\X��ˉ.��c��!ry����s�n�>�C��7�b.��PN�A;6����8����m��#J+dR6FG�p��3�n�:dF�a���O�U�<ۦN)A�e�h5h�jH�� ����,���`��a�gg�l���9$F
vn�F��8Xh����aj����"r�h1�<&�Y�fE"�9�Q!���G��U9���}l?���j���3v�W�V@?G�^K+��?�w�ۥ�G�<u�U|玽���I,��D1����ӎU�6S@����U%l]S��q�c�VP��E���"����n�P<�Lb�G����v:�.i�+�_DJ<� R�(DnZ��#:�.�Q
庅}Se�+]Tz�"ŊtO��*)!����˄��<�����~�>W& ,��6������3�"c�Rng<�v��!�X����A�������������R$Y���AV���[����\p�6|�;7��
����	@tȞ� ���HЫ/�O�x�Ӟ�W��r�f:<�/��?�ڛnG7��C�-�c��b+-.g����\�m��ٿ+)�_��7q����@��Jj�ЯNM�ͯ�h�*	L���IXS���4��ʧŝ�?!�0D����/@'��.��� DhM��mZ��Т�^π���X����nل��ދ�s��Ԟ#���5��=Gk�_����W�G������1\,�c�>�T�u=�o�Wjr�i�%h�B'dq�jwu�w�H8C���`�@:(�|<��O����٫�T��݇�H���i\��o����pr����r)�9qk.�c����u/Ã�\M	�`�*c��Q늾��+��|調�5?�����F�ل�s��F���L�%vВ�"\JQq� ��@!m*�dM|��ހ��[o	(�{�>��p��)��k�
َ�K�%<Sm�6�w��q��0�H
'��RAӨ"�j��i(��愃�-��m�	Dv�GB
�~&sub�A]��\&�t:���'���/� �y/�'�C>�j�e$/�P�?�e�9l;}3�ܺ������h��o�0sH1L�������\G!�[�ڱ�r܀��!��e��<�}{�<_�$5q�^����ʍ�m�q�a��pr���Z�6�g�m����4	 �I��.T�7m=��z"��L#��;g�����������,��ob�.���*/}��jn�}ϩ	' �޹?92/ �ZZ]�jFa[wR#�a-Î;�J��:��%���8q�.����B�1�򙫑 $M��r�b�E)_����	԰�#�Q�n7�ͤ��D;v��4��V��x���3mL�v�G��n
`�n�I
�x=��a�4� J��u��E�B�#:<�0�/�I�6;�M���9�x.��at��ۗg�o�:������cL�,��:|vz��-`�?����Q*�J޴\�~Q�p�|R�-� BJ�m#ɗ$�� ��ˠgz�E.�-ńL@�}Y��a<X;-n���H�HE�[�s"4����LMH�%��⑅%iX�H�gs^�������(�K@��I��)B�p)f� �6��n��¶	(SƉ#�/
��=<kҎ��c�MW�/{�f㮣U��u���Ѭ�ۦ��� B/�j�?��iJ�s'1Z��͛�g�8p�8���5�34B�i��љ������j7�������X=Q��/~y��x�F�W��;�4$8wͨq�;���ql�J(/6��ʾ�]��P�9�U#|�C����JƎ�bw��l��%�{f����80]E�Ќm��VA Nd�;:{��*A:Y+i Hʼ%z�~?�.iKk��x�[^���6&.i�c�Le�������7T�zl���H��VY�#��`V$!�0��c2['	�\	�����~}#�0�`Z����Rgn����!�͢Ѩ���ʵ�s���Z-�{�<�h�FbM��N�ψ1�1�iU	��1�5��FKL3��}�`պ�[�v68>*�E�8��Q�o������*���\s�6�ru�ۮkÀ$ �zݦܓh��2�g�o����B�*�^�h�L��<��:H�d=Ʊj�gQi[Jځ�F��;���eÃ���ۼ���3�W<��X?��nG�Jpу�+Y���ric�V�W�Kϯh!��恱�'���jq��� 4q���uw��'*X�S�vbt�m�Rd��kM���p#ͷ�1)<�-kF���5�5��<f+F&eHA�D���YP��N~�PpB��sణ%}�.:�xPL�5|�F!;~��\���Z��/�RO�	(Ve����PLj�]��1y�{� �3��g��y�*��ˤQ����||�F�0�Ia|lD��CG���w��@�t	?���{LB�� c}�X1�NM&+!-R�'1>�@�b�@I�9M� "N7D'��΄"��W�)�ڤ���Nb���lD&M��s���	�"݌�,2����n�T�:�\�Y�1}�vu����x���]y#�V��L�2��h�b�)�l��ߊE��	��$9]�s�=�9���'r駯Rc�L[VH�&r��#|������<�4�~(m|wǴ���]��b]�D!,�]l۸�l݈s�9��<j]�#��|���H�7�>����H:��LN@*�?��"������.؊|
h,�ż@Ť)lN7k��3���{8#_@ϲrZ�y�t�s\d�����a�71���mǱ����;��/��-X�,v"��M8����(`����y	���jէ
GK�Fn�=e),/���?z�|����\S<n�B	������M������PAK�MyI�׀��Fp�	�hءG,��7q�!�a����� \[	��]9�\;��fB�Z��e��ҍ͵=	/�N�r���B6_D�n9������(R��`�`c8i��9��9��]���ah��UkW�0� �fs�vB4[]P���:it���1��Ait�XW�k��t�V�Թ1Z#Sߘ!���F�Ӟ��<,��L�B�V���q����],�;p��Tq⢗�hG6��ÉF,Y-�-�A슶��{-��a,`�Iy� �
�^�{i�i����{2N���������/X�������X����`ї>������bW��N�:��)�djV H�!d�$k]@D�r���5!;Ќ�16�aY)���2��O"���+0��#t�1��cJ�ņt�K����\�Nm$N
-xH���>��Vpd����(7zH��[��D%Z,-�'rҥ�o!WȣX,����N�����Hc��#ֺ"�&e�E�s��iVfa��9�?�p���ga[���`�ty��C��Dt�`gI����R,b��[���/�|��0  2�`p7��_��c���΄P.d��=Q�0X�FB "�,~��V�B���a)J��BdΊwL�,*i.��?��
��cn�PcXP��%�����x���������%BiI��o�|��Z_�q�\�� '1`�I�zʈ1�uq�C�ċ��d��|����g�(G겧�f~��8�gf�N��>�2<����vy
.A&�5��w��]�(*
�-m3xЃey�6Z.�ۨ@��XQ��K�A��3���@�=��,�)`���������� ��B�����6jH1�Җ���m�~6��p�δ�����F
�ܵ���װ�dI���F��?�@�m �1b�L�lN��6{}������M�)@���I~��p���޹�J� �����x����* $vs��4t�%�#����a����VֆP�H/�h���	�o��_�/3�E1uJq�h�E��	j��y\ɮ?�[Е�UK[�=�^J7T����)ǆ�r�&riy���k�1�؝����I�3zX�b��E�۰7o����;���2�E��
�.<4��0�)������kve�y��<���LXð�'��>P��2��Ihc�E�ӥ��⮻�>qR�1���"l��X��i��tq���\GI�|=��Bm�+��6e�%@�y�(3    IDAT���_��#22٬���Q3�˟�����[F�5qΙۖj����|i���+�t��������W�"���i$@�;1n�w7�=�r��UH(�(�>o��n����찓��wX��`V��pᶕ�c�y@И��hV��b�@&��6a��kM }�E���1ۗ�)V&">x]��C/Lc��`���8�PC�ݓ)@Dj'%��0H�a�N�Ģ�	�)����x��ɏ׾@��$Bu��Yҹg��A���
V��De���ۑ2D	C�BR���nQ� @j��m��gsB�Q_o��>UIF
:Ka�M<�ۡS��\~R�"�$��X �`@����T4�&bF}�S��B�i�QR��*x�'�&o)#���/t6Huc�e²9U
�ޘ�i+-Aзc�9�j ��(�'%��U�ժ��ɏi�LzhM�xBɡ.�>{gm������RL�7l*e��_�6���ta�\c�a<�Oƣ/X�-%�Aw�U��c����9�x��0�,�e� F'
�"sc�&�X�O~�E��g<��_�^�
�T"R��4���P��}�FG��d���s����[�9��`qz3����$֥c�9uښ1cr��"��B��}�o���4�f`�ы�z�]%p	GM�E�̕#�$�������R�d��	�Jddt�?y3��]�B�]Pw�܏�|��{�#;�&4=2	Z��"|J���u��bH�'~���Ӷe�џd��˵ ���'e��iZ�KLx�-!Z���	�t�h���*Rq4p���nU�θ|x���Gm�S6�ƪ���B]4�C�U��锁�R[�n�����q�39�-�9$t�J��W��׀�@��}>�A�^E��q�{(�w]��9M=��) �`Dn;����\.��v~~�� �#G��iG�Ӆ�ɣ*q��C7���r����tG�j������D6[B�ڒ�eL[667B��sc�!B:��B�� $��]~)�X5�]M��9{	����K��@Y�% �@9�K��+[�;��St j�"��j��[N�;�LH���@�c!���u7���ؒ A��V]
ء���+
/8X^�`4��5B���{��H��)�
_��ɗB��4�ahXH>ls�.j5`��,N�,��+�@���w�M�R�� =�ۅ�L&#�j����"�f����"?�/�Ϥ�0 k"p徒��C2���>)�:��c�2� h���F��|kѧ�Ќ���w���44N��/��! o)V�JNm�o�b�R���㾋kdȄ��X��pd� ��� -
�E�	�:0P�P�l�Xh��n��~ ����x�$D)�s�d"����i�A읚���",L�)?I@
�5� v�E��N1	f�I�vhl`8�Cu�(����wbӪaؤ#�16������+��9�G<�b<����p����4�8p�,�!#W�T����u��җ*"Q�(Ԧ1�cNEmCi�{����g<C#�@�٤��T�����_}
���&��#��R�!�	���v�i`8�F

�'fp�����ϾØ�)+v:~3�#�S�����o^wZ��<4��3�΃��"�H�OJM\�ө�r�o����s<�Ŕ����:<��U�&����w�Ƨ>��}�q�&6`���RzC�d:��j&��~'_w���B9V<f�,C$5-�L4����mA�"͉I�q_�n��8]�7RF�����)�霞0�����T�R��B�d�A<������
X5��u�^@�]D�*�DF���ec&��N�-[7��Pqi������:�e��9��p�w`r�ꍪ�k&�C�6���RI\�8��5J�b9�d���>)��t��}��+^����L����XBK[=����Gfw�< ��2dJ$��eŪXB()3l�N���m&�29	������P�Fь����m�Ga4�s�����K��XZ�_~�.�_~͖~��?ޱGq�Ћ#q��oE�n��p�QT�<Z'�:��u�>"��&��,Z��ǲ0�i��������a�"�B�F!cb���bW�;�n�`T���а��8q�v/��P�V�82��L����>�9!����75}퀀n''X���(�{)�����.��Be��ȥ���]�S�)�Y(X&'�kJ���鍞d��˴�A�a�e9�rA�t��BӲ��焄�%�[�<˄��&f�p�uN(�E��a�D��T8���P��W�������O���B���T�����O�����\�5-*f�������k2X�~�9p���K��;�o���k��C�e�=Ǡ�<�Hsx�C���]�&��\Ymӂ�Ʌ�Z7�5�{jӰ����jmIg�L�یK�i�?|�{�No�E�L���my^	r)����������a��A���y�Ö��������H��$��)-ɣ��_fΰ+�"�tZ�]�����~)�^�����C'�)�Q6�Xv�9���O����Xl��/C�j�A�*}N�5F)��c�w��Z&�"�p�.y�Y��;��f�0�MO+�׏�ѫ��?��XL�i����9�`���C!�AS�d�t�B�W,�y��u Ǔ�u�����^�|}���E4Aӽ����k���ny�Dr����5<����Lzp�#0B�S�8��<��2M=���	�����?v"�?Я���6TP
��1ilp;H�#͉S�t:+���|L��Z_Գpz�i�9)c�N?'&&��)��g$0� d�����)�>4�JK��?�|,�'��iJ&)�aD���n���FPÛ	�=�W��8������,Ⱥ	���g\�p���,<��%��Xڽ_�
,�_��.���s~|�^>�E\L���|��s7�A�)�I
V����B�F)Ĩ���!�E���4B
���ݞ�ڛ1Ƈ��.�|�B� ri�%�p�b�.6�^� D/���j 2��Znf�-y�����9�l]�jz�Б�q�a�U�]��th]�:��U��;�@|mڰ�3�9�Ky��g�s'�~�T�O"�&�I\�t�W�}�A �]��c�!����L��'�.��%K�������T�[O`4ʢ��?��d�!Z�5��+=�|�����2�� P�˕\:�NOW���d��(���1c�o}����)��4����¥�\+�`ȷ�zÊa���������:j��ol+���G!��H�<҅q4͢��4�K#�v�y�8������q��ʸ&6��g�z,Py�ո���g���z������!ב�i�ׁ�a?���:x£�����p�J��=��8eܺr�19;�((�tp�X��;�S��z�����{7�X�,���`N`��v�a�33aN$8��1br����"l��K�x�ˍÍ���l�a�ox�U�s_�F,�DOaz��!�P�C���}'59�G��(�Y�n��:A�z!x�\7�9��^�9�!<��R���ɴ��ў�	��i�d'1�}y`�A M���S�p��"�`�F��TQAB�P�ރT)�J'��Ҥ��;RC�t���$�N		�����r����;g�;�s�\�#_��Ai�+����:Ł��&�g�p��3���L$]�-+��M;�#�W�^�m\�;���-x�8��%ѿid�t�4�K����ی��'7t 5�;[��XȄo]�����
	<�y)nx��Op� ㅬ��|!��(1(��h5�-P�}K;GV��)%�Ko}{��V+|��������n�3Z���#�6�pT��3P���q0�L1X�����+y\�\E��Pۇ�=w��'�4�+�l�߽�+�����,��M�xAPzA�珴#VΒ$Yhb�M�����§�ץ��י�&~m}�}d.�b�'!*8LKRx��݈�[�j�_b'#�~�+V���;�����*� '���u�U3ٵ�J ,�ӥQ~~bU/�-�-�y�����?0�)RT8���3�=��B˭cy�ɛ���&z;��-7M|�e&.��ٵ��j�I�K���f��(p��<���4�M�0��s�O��./>ʱ����n�fG6=����XJ3Ns��~�jӥ����B�7��b�:nw~�۽��7Ô@�k��RT� X�@��0�LI0�>��Ұ�3#}��[Du,��lhK&�����[�m�.՟d�a�<؎[���J�uN��͚�D�K${�n���Q2i�q���@d�6�=_��{�?M?�/���q]��BN?�����3�}׿ag��=�r��M���V�S�n�y�m�C��b���bBX����@�aN��.��n��(8:��ڸ��L��R���!���%��z��l���� �3��k7���8ȹb�\|7�VhWR�𽝙��>�ISs#Μ���8�7%G�0V��-��S�
Bt��+筟�Bϵ���r	}g��[�]"鵹hcT��k%���봨���R�m`�VY�5N��j�a�FІ5���$��x`6��DW�[�y�t��,HfM�,� ��
�!�vo�P6�ɂ�Iq#�|���X,(Lb�C �%F$S2���j�þuϾ������<�k+4���t��m�-����E���k'V|���j��U��js��-c�vY�F<?QD2X����b+���L�>VO�At�`�j�)�-�7�1��5�Ag�����$�%�X�Fe����Ej�О��Wj+w�Q����$$s�E�\_c���:��w�HXZ���B����/-�*%���޿{�eX	��x���x� c�V&y{��nlQ=QRK\���UYX,,��w��G �'eGG��E]X�J���2��\?���F�Fu���n�u�Q\�J��Z�Y�*�iSPy�l��D�q�P�?��7I���ْMV/�U �L��A\�*�aW4�0ɼ�����0�_r3�T���/T��A��?� �8Z>U-@��&��(`�7����ZR�c��(�h��[���D��d<q���ͦ�{��KS�8
�0�"&[�v��]
��}SXaQu�9���A��i�jN�����j�p`�"�vђW��3�R�:G9m�|q����V��������vџm�̓�5���Tx�ϭbn���C��ߨ)�������
p��OM���/��K[�bC!�5�aӜ~E��<��#ն��7�UW�Y����5x�)ӵ���3�K'�䴒�
����A�
$\�d��+��<	� �`�~W�������F�'A��z�u~�a�-���`c��)@?�g�$�｛�G�~E� >>�7��p��F�)�RE���+)�ފխ�E����'�W�t�
z���۶ʠ�G�d�����'k�-J����p��(��w��[���4?�fR�t"�ҟW��~�H*zi��r�{�Tt���rO��RO��}����)4'��A@�v�.�����;ȳ?N>�>�|j���	�7[u��fg�i4a�HJ��Ӄ4�9v��陔$||f=��wݍ��M����B��s_���"�,˪;�UZ���1� d}�wK��ON�'� ��-��r~�s����1.ϧ�g���R��C���n�����|v�x?�
~,���e^�1�{G6��Nu�~�G՛�wFS����c]Z^��9�)�I0W�W���wI6Dux��3�m#��b�A)4�W
T��"�-/���<����G�>�ǥ四��q9�n���21����o��l�����ޮ�Ϋ䃦>�q�V��=�t�c�,�/�k�v���)*B���As�%H��']�\YT
��J��QR��A�M����ؒ<��q|�'���+d| ��2���r�4˻��X��\�`����s�����c�h5�+%|���ZI&�";�O�U"V�}6��S��_jɯ&�6[W )Y�ِ#o�.ۢ�`�1�Qa*l_�|��j >;@�Z�*>��<���P�i_����E4;�轌Kl�s�ί���bЫ\��zq���VTн�*؏9]�J�7�����B��,k�f��l�n�_�v\��\]1���}�%W���Ħ��vA|�c�ږV/,N=d��8�G��**��X������f��򝁉�)�����Kw�\���p���2O����kD�Gk�Y>�o*-�W�RV���q!1�RU4eδ�J�cso%<�3:�0�u����Ԫѳ�Ф����v_�S��$�ԣ���f�0�x����.X��
_"ڸl�;���(��'�ѽ�b�}8�"��s�~�Y�PƷicL^88��6���$r-k�=�� ���~�vp�T���m���@��nڡ�XI��m���a�Edv�散ZV�yH��>�	�'���/~���f|l��Dd�*a�J(����{]��w@�H��_^�~�ׂ<��|ǩ�諸�w��q<�j��K.�{�53�"�XVT@����5��N�N�0��v�N��Ո�#�)T�4�_;�<w����5�sf.���qĆ�1mfX�I]�3prQ+}��]�s�,d'%@����y��v=>��ѥ��.1���77Е��5��O϶��q9H		nĘg7D?~!��.�c�p;�����&������^5Qz"\�ߗ�@߫.�%Z:��K����n61\|�
��BYD=��F*&Ɵe�+�CDEd���=�����U&e���PkdW)��o�[ؑԛ1��rNp��i��W�ƣ������u��#��w�,�j<�b4�����'P&p��]����+��ޤ���>U�8�^�ᷥ4��0��RCk��6��?�>��~�9m��� Z��`,��M�T�AZp��4ɽ���t�[��I� �3�F6��ϧU0�n)� ����܊�'���jH���a�R%e��^�^�[2%���a�zJa�%�����S=G<?X �̈��ƚz}�έU�)�d�&\gtx"�P
I� ц?�A�S9�.��^��]4���"�����#	��ƈ6���_fz��nyoL}<��oͺ�ȹ�ۏ�m�"�/[�`�\;�������\&Z}�8d����?_b�k���Hu��B� 1��e'A����z�<�Bg�4B�׉�|TЯ�&���qL��7$.U�;����{Ŵ�8�`@�q��!������&C�\��I������F���9s�m�|4H�ӟk��̙�$�s�}�7�6W[�
��?���t�N_!Mw��:]�6�x�h1�{��.d�^���qC�Lkz��� �|�q9zqD���� v�PE YMwX��_7��u�����E��@�-^B�:rO���֎�6����N\G��eE�3B�ZC��9�tF� S���)_��p�����V'�+)�� N�sh7�m�N�~�=<mmnAh�_Kb�`�qk����qM���	��W0�3�#���k{t��{�[mt��nrtE�c֓��Q�6촕0q~�I=DH�v{���ޔ~9�1���a{<q4��kv�!`�5�S~����8����s<ݙ�h�(��������Рr����hp�l7�̡]�?nR�U[���s�nXpՂ���Y�P�[�"h�5D������̣�����I�E��,{�j��Hl�ۧ�FRN�b)r�ߑ{��ܸ8�iЍ��R���/S�L���+Sq��=+���q?�ze�H����^O��*�#K��C�:�������J�eWi�Ɓ֫�)�:ڷVrC�H 0Q?7�Ǡᴥ��5�ߔ2*�+Iu[[��M�Z_���6,6�Ҭ��H	�F)j9{0s�S�yp�;���L�nw0�_�4�eL�Q�h�!�3���@. ��Y��$�a��赳�ڍ��M�w�m������"wռ�\��3�)I<����Ғʜ[:;�G�`(oC$~�ȁL�s鬘�<����J���燡�c hp�q���ߩҿ�rq�f5B�e��S�l-����+|O�'�v��P��}��]5�d܀�A��f����T#��g=��o��6`71>Ȩ��M�ʾ=���5��:�P��ث��Vw7�ª��UG~|^��e;�q9 H��%W ���_�r笷���9ͩ��b �lZ����w���)6*+S�y�
���D��L�����u&�:��WUz�ڮ�5�����ٺj��QS��v�N���֢W�eh� ^k#����I[��g�44�!��`�x�Q�1 �[k]J��ӭ����2�r����~��K0��Dky��H����޵m�j,9��@����폄��3;I�0��i8��|j]ꇡo;���2�(i�)]*�A�0?���]tt�9y���BX.1�u� OZ����:����Q���]����A��T�U,�\���%1؜r�dTcH4w�Z������,>L.�ї	�-��KT`▇�s�=呱�r���/߽hM�<���H8�gj����s�z>B��^� m#wcm:l�@�YQP������Ċ�n�='�I}:ŀp�9�q��l���js�Gu����'������jo��:�����%#�k&��&{j�)ɍ��a%���^�꘺нM�8�9���1���8\Œ׬����.ivPÛ�䆚�>�e�
�7��nq�B6f$>̂���'�.�Yd��ug������q#$60���7|c���h\�>z��}H=��ڰ�c�ZDz�B�ctJᙐ���w*�/�.�Vɩ�(��=k���ѷrK�(�^�3�h�;7!ۋ�L�`��0aݯ����M-�+�F��B��<f�����z�M޴�;䜨@�-�^mpgD���9~�|���ha��_,*��/�*ד������\��g�_�yꕚ��l�y�"�z(��63�|��M�B�X��S�Ƈ���[��Й!��.�F�$Y[��O��&_Et��$��{��Zc���O.��';ڊ�B��G��j��j�M�5sf��.��	�:L��(}�S�İ��Gբ��2�A��Q��r���^���@Ud�Q �����x��}w��OO"U(�e��$��F�e�CN*1�@ZP]Z��uy��GS��TQ�\��vӕ4�s�:��D�ǩ$s���_P+pf�����k<���
JT���Z�~FxVL�Ӹ	&[c���H� ���w8s�ΰ��Sz���b�>�,����nO]x!�&lUg|�q_�I���w�G�q�]"k�*����]��
����}W̋�H�;n���m3gk���7Nn���N�V��k���g��2�}�~x��*�,w��}M=�&!��/3��I�D3�;%��c��q	�w�m��|����(?���},��;��G���2�����u�"ヂ����qk|�^�.���M�X�O��R�N��*��)w+I�'*��IK�R5Dr���~�[�)��@��D����rz�nMY�}'�ph�!G'"{���x�v�8a���T�dd�o�t���.`��1��;G�8!JLM��<y��}8*T6R�j@�T	���Y���E���e'6�6��is��Wcn[�"]�~�Mƙ�8�'U�K7���m�{��'n�JN�P�[��J}cj���b�.�{Ê���!����������sP�X!�pGO��4�$�]��nϟ9)U:�2{s".� +茲�7�A
�ܩt��I�橏���7���s%����1l��g�Br�>��h�%�D���k��;=�`E�6�O���9k>S��H�~�� �a@U�Zg�Cjj��3x�����u@Ӽd.��3��x����@����# ���y��s�ٔ�}�J�'���}ۅ����O�l��T�	�Ի=�L�h
l������Ӽ&��?��vk\'5}�`Q�����zK�G��pۀ`ll�'ާ!s�@r/}�sZ�ߔ��w��Ti�8g�rm�����W�?(��=��_���k,U���V|~�rMa�W��|`O/?cp-A$(YyzE
�^��2��ñ�Uq_���Z���i5��":<x;y�)~q�X�P�#�O ,W"�;����U�u�"��e���h�h�	�9��W9�S��JyV1��|����Y�D���,\��VtH�A,�O�i�����d*Z`߲�����>��Kv��]Ƀ�
��v�f�I�~j��7�q�_���~i�0l%w�ʾ��l��78�+I�43I����Y1��t��&~��c�f���a������ p��r��$�y��A1ش�
9�	m�H\7Ë�?��љ��-f��(ya���;J�����☖� 'v��:eM=h���N�"�qC��1�+��F\�:����M�ӆ��+,������k+�s,�_7�l�����R��sl���=��p��B0-�.��B	s������o�*�Iؙ5D�o�O�+��=^��\��Rzn���Q����xq������hB�\���y]��K�<���2���R�Ԡ���/�_ҿ�I���%�K���/��!��Ӂ�s,_TEU���@�����,C�PK   *��VJ�1��  >     jsons/user_defined.json��0�e�k!-����ɲ�MsQn�d1�rk���.����A��6�+�K����P����}��u���f*ׅ���Pu��6��]+M����~9\~����wyw�1�P$�V=����=�o�q;A:��<M9SB:9%�C9�N���Ʉ�8ϸ�� ����:m�N�z~�Y�=�:ם���[��W�bQ�%�P�=E��v�~^���\�)�P���.�O{�>��8GW���P,�M[k���������K���3`9���q����F7�B~+k込�f�>���8��/��<�5���WѠ������?����~4���g����g������߷�g���Y��U����=��)�k��GX��Jխ>�E�eY������̇�C�R��\r�1��"uh��3�O�0dD��y�G���)�ا��+�'���	�����'4tC�I`��M<�ߍ�O��oĔa���Mv#b����0�0t,�6�����o���O���=�PK
   *��VX�EfO  X�                  cirkitFile.jsonPK
   ��V�4!V��  �  /             DO  images/1efc6cd5-4b9b-47ac-a031-8851919f3fa8.pngPK
   �}�V�Uˮ�# s5 /              images/fbb65e9c-f417-460c-abe8-d9c00fd6ec79.pngPK
   *��VJ�1��  >               16 jsons/user_defined.jsonPK      <  ^8   